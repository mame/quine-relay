module QR;initial begin $write("%s",("let s=(\"Module QR\\n\")\nput=s\nprint\nlet s=(\"Sub Main()\\n\")\nput=s\nprint\nlet s=(\"Dim c,n:Dim s As Object=System.Console.OpenStandardOutput():Dim t()As Short={26,34,86,127,148,158,200}:For Each d in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import :wasi_snapshot_preview1: :fd_write: (func(param i32 i32 i32 i32)(result i32)))(memory(export :memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export :_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(d):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(6"));
$write("%s",("21635.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n=(c>124)*(8*c-40146):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^"));
$write("%s",("nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^6"));
$write("%s",("3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3ciaqp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]13nfa3(f\\\"\\\",2):f(\\\"\\\"{#w3nga7(f\\\"\\\",2):f(\\\"\\\"{#.x3nga51(f\\\"\\\",2):f(\\\"\\\"{##4nM3sca3643qw3yf6dx3kca\\\"\\\",2):f(\\\"\\\"};l4tda,43z3sma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\""));
$write("%s",(",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCc4tC3pka721(f\\\"\\\",2):f(\\\"\\\"{#DNE;34da. A\\\"\\\",2):f(\\\"\\\"{47eaPOTS|48\\\"\\\",2):f(\\\"\\\"{45oaRQ margorp dneF34baS^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'46%8-ca83737ba&J4-93bgaS POOLv87ba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'83[83ida&,)-96ga. TNUO655fa(rahcX6.%4dgaB OD 0096ca&,\\\"\\\",2):f(\\\"\\\"{83ca)AW87R86qaEUNITNOC  "));
$write("%s",("    01)66~67D5/n>deaRC .>34ka,1=I 01 OD[@8caPU?35)83va;TIUQ;)s(maertSesolC;XHeN3$ra598(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})420:41pa9191(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})84022HxX5qca69mIy[Grca08<H3ea5526~A[83odamifR4.fa93623R4[83nbatN45%a315133A71/129@31916G21661421553/Y35wa%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})867\\\"\\\",2):f(\\\"\\\"{3ahaj:+1 j@a45baw:35935baW:35ba\\\"\\\",2):f(\\\"\\\"{:35va)(esolc.z;)][etyb sa):9[83;ea9746(?au4[83jba,t4[83jea!\\\"\\\",2):f(\\\"\\\"})8j3aca~~#4[83jea(rt.w4[83jba)<5eda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};m3ffa~~dnep3ira~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a73k$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||23kda#-<r3kda||i+3nhaBUS1,ODw4rka)3/4%%%%i(S4c~5l[4yPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(ev"));
$write("%s",("om(dro=:t elihw?s;)s*:5pm5ww3kn7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/GKa|atnirP/oi/avaj lautrivekovniJ3d/4k[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);80022<i;(rof;n)rahc(+L4s[2k+3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'oa=]n[c);621<n++t4aqa0=q,0=n,0=i tni;O3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'kc6awi4asdRbQeLlxfvfElRf<bedRb;fPD;agb-a|dzdxdRfGb8aqeRdYd5azp4i;agb-epb>a8adeaj>aJaRaAdteFbaeIfOa5aac2gL\\\"\\\",2):f(\\\"\\\"{6f9ak+4aLa7a;a4a<aNhUmkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9ak+5d6cRbC3gYc-f/aof0fRfCa>a5arm.b2e6aRa;dp<ogX6Eh;aTapc4aLcEewiof6amc<byg-f3msbuh|b*bWfybxcxc>aGaUeAa2a6a\\\"\\\",2):f(\\\"\\\"}g7a6a@a\\\"\\\",2):f(\\\"\\\"{g:a?aMbKaKa6a?e:aS72a|gZfMbbgji>a:b1a-gSmUf\\\"\\\",2):f(\\\"\\\"{bHa4atc2ij8KjVLwbEc3b\\\"\\\",2):f(\\\"\\\"}bJaMa\\\"\\\",2):f(\\\"\\\"}bJaD\\\"\\\",2):f(\\\"\\\"{VrJaJaB9JaMdJa8bTaNa;a8bErKa8bEr8bTaKjPtOa:.j89bKa-=hJTa8b=.Er8bj8\\\"\\\",2):f(\\\"\\\"}4JaLaJa8b=.j8j4eoa8bNa-?j8:b+bVL*4aiaKNJaHaJa;3c/aHaJaFdTB;a-=Ua:aUa:aTaNatiSfQf;m4a.|sbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\""));
$write("%s",("\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'matiDa-a|bn+-aB6asaYYUe>atl\\\"\\\",2):f(\\\"\\\"{gKaKa|gZf$6cgaag2kkg(6esasbuh*b-a/bxcHa|f1le3c4c\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{goh\\\"\\\",2):f(\\\"\\\"{gvg1a-g\\\"\\\",2):f(\\\"\\\"{bHa1lRf-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?a\\\"\\\",2):f(\\\"\\\"{gJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1a-g/bHa1lxcpb7anb2b:b\\\"\\\",2):f(\\\"\\\"{g2fuk@d-aIfAkxcHalgjghgJk-aUf/bHaviRf-f-gSf|f1lzeSgviHazl;a/aBh<b*hUh<apb/aBhUhnb<a.H:b\\\"\\\",2):f(\\\"\\\"{g/aBh-f-g+gH>Ga|b1aji3b:b\\\"\\\",2):f(\\\"\\\"{g7hHa1lHaUeH>Ce|bxc3b0a:b\\\"\\\",2):f(\\\"\\\"{gIa|bzeJa|g5buaQbvi<b=a-ahl*c3bxdUem3aea|b9ai3era2bMa7apbphnhlhjh9k3fAaAdiFPcgfvfMhHh7aEa|bqlolMahl*cEc,dJa>a2aIf@jMgMahl|b\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}i+cZh6a13iWa|b\\\"\\\",2):f(\\\"\\\"}iFwgX8g/aBh=aniRa2uCd2ukb.B\\\"\\\",2):f(\\\"\\\"}xnink6a7b:lRfwbCjUe2bAdamGF-bhcQplklkVp0c/bxd;a:h5j)?aea6a2bP>emc-C\\\"\\\",2):f(\\\"\\\"}U6aoo2a5adk<O\\\"\\\",2):f(\\\"\\\"}gChvmdulk6aSh|mHa:exl8l;aPlQa0/Rf;M<b3bxd6aGh\\\"\\\",2):f(\\\"\\\"}l5ahj?UiivfYgacPa;axjccUIpbubldic+d,bnbpg;j9jEc,dxlGk;ktm<b<b<b\\\"\\\",2):f(\\\"\\\"{k:bqk<b<b,c,k\\\"\\\",2):f(\\\"\\\"}k7b-b,kVvSg3bDdilnj9a7b6g-a5bs\\\"\\\",2):f(\\\"\\\"},c,k=a9a7bubxbs3ekawSkl,c,kAa13ceaQD8fA3c/3ifaJb7bd%3dkaxkALCk9a1Z^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3cmaiiXk6j|l,c,ki3a3a-a+bhh.bfh,c,ksbHa\\\"\\\",2):f(\\\"\\\"}gQk@lkg>l8kykEa3a6a"));
$write("%s",("nkum7lmji3aiaNkgl<bzeACc73ggasl3a6ab6cka;M7eYjXiVj^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3grb,lmj6a<bii\\\"\\\",2):f(\\\"\\\"}j-C0G0S9K2a2a;MAkzlHawbCjRf59nc:e7b5aWf=aKcFVbl5a,bJa6a-bJaJaub7h5aUgwbCjHa:e-b9a9b9aslAkyg>am3awa@a@aAkyg59:a|b9a0b9a59VBa?a>e|bPg9bJa0bAkyg-b9asl9aCaAaJa9bAknbJa6a|b5a,bRf:e-bql?6-ah<a(aik0G0Sti;Myg8bAdEh-a;M*b.bbb-a;Myg7u3j53acaxmf6crbBkrmWjpm;MKc+i3Cxd6a-b9a8b9a7bJcJaybxnu@>aJa*c@dxc?b,bYI>aJa-b2mteUe59<a2b5aDcR0:atcJaub5aEcR0?aGF-bVgRfn8aga5lmdJhm3akaNkq?0G0S0c.4as3awe<l3apb;awbCjWlbkyW\\\"\\\",2):f(\\\"\\\"}UwW8Ix4Tp<Oa-x4|U6/QmYl3nco-mtnro-aioN4co@mL\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"}?GrIcbik0GxYd=vYN+d6sWdUvwv>yK|FDaBa|F7va@,t1z\\\"\\\",2):f(\\\"\\\"{8Ea|bErDq\\\"\\\",2):f(\\\"\\\"{Bjbqp*.a\\\"\\\",2):f(\\\"\\\"{9oz\\\"\\\",2):f(\\\"\\\"}KDCU9oE:3bj0;rA36sHoeV,b/I5I=CAp4IZolRPaDaib@aR6rpkdt0I0QAjbvb9B=aL\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}C5p@a\\\"\\\",2):f(\\\"\\\"{/1t,drqHqDa|OYaEa251bDa2b=atb,t|btSj*48=5v9ab@pnEO|6Y?Gtb;-Cymb?GnrC-n3tvAav\\\"\\\",2):f(\\\"\\\"}H+fvqK??l=S4QX8|7b?Ivr7q88dwUWsEz,P=ab.b+i2\\\"\\\",2):f(\\\"\\\"{@ae5puTapthpubgT3b\\\"\\\",2):f(\\\"\\\"{q/=/|Ea|.QDub4HP,Y;NT*6e$dTaiuU5,@COsl\\\"\\\",2):f(\\\"\\\"}7Gq6qlbk\\\"\\\",2):f(\\\"\\\"}j8h+VN6l2I>aC6u6Fawt<a-AmbJoYaLl@tQ0x+gttbnD\\\"\\\",2):f(\\\"\\\"{bktu<WaZ\\\"\\\",2):f(\\\"\\\"{9z\\\"\\\",2):f(\\\"\\\"}HbM2*7,n@xbYp1:-i8+=u*LGp6s1-X-=uSajbA0<-0:Ny2blbvbk2Fa1t1bRaE?G5CpA\\\"\\\",2):f(\\\"\\\"}fbBwDa+b6rDS*b64W+ttRGbbabDCtU+u0s\\\"\\\",2):f(\\\"\\\"{*BaYG15T\\\"\\\",2):f(\\\"\\\"}r1Wt"));
$write("%s",(";;cXMLYtW5Facb|DRa6wybUHf4v>PQLu,l9p1b2bPUNa2<SxSxt.N>RG0szzh2ybBaQIi-QD.3-qA1iQ9W+WMD.bU3Nou\\\"\\\",2):f(\\\"\\\"{ac,6eEckb=rGhEagbr.\\\"\\\",2):f(\\\"\\\"{8\\\"\\\",2):f(\\\"\\\"}buydb+bAarpcUaUCaYaQv,b:t70VxgxY7HrEappP=U|Z4;.u@QJjvFa;.?G36iihPopjbxL@albau9J\\\"\\\",2):f(\\\"\\\"}WuB\\\"\\\",2):f(\\\"\\\"}bD|Falb9oPq>wDaK5VaH<sqD1r.k\\\"\\\",2):f(\\\"\\\"}S00\\\"\\\",2):f(\\\"\\\"{KpI:1bJCkhWap/djjbvbXxI,d+kUiiH1sSOoS/DaL+AqWo?GYEVSvvjbVaRSdjgqkqLSF\\\"\\\",2):f(\\\"\\\"}ISIo\\\"\\\",2):f(\\\"\\\"{?W/7oBpOSDaBr9bEao1jb-nUt6bCaNaq3a8aDBUamwr.NO2b-SVa,b.8BpEaDaLsGaQ*wS|O\\\"\\\",2):f(\\\"\\\"},sS.8jvDqs-jb9Y9fOaVa+bYxBpEap1|4=qXa-\\\"\\\",2):f(\\\"\\\"{?Glb,q0wr.f\\\"\\\",2):f(\\\"\\\"}r.g*Io|FW/Ea>jTaFa4bSajbQaW+xnkbErDqFt?G9bf4a/aiv;jBaEa5bIo97s:0AW/EasYN\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{b6rO,0=Pa7\\\"\\\",2):f(\\\"\\\"{J-QLs5aYb*RQLubDaIrHo:BjbDaswBaEa:Bjb1"));
$write("%s",("rAa\\\"\\\",2):f(\\\"\\\"}xQLub1rEa1bgboRX5lRF2Ea\\\"\\\",2):f(\\\"\\\"}6gReR6bwbDa7b?nwvEaXv.bgDt>tbVQoKLja?7bF,Da;pZaqqX0ALjbD82>Jnkbt0OzE?aHBa\\\"\\\",2):f(\\\"\\\"}Qg<4JyQ\\\"\\\",2):f(\\\"\\\"}pnx|b9T-hkbXynpYh0NPoZVX7w?ibx32Z@f+ciblvhbmbzC+-j65w=aAL4b|K7rc1,b<at0ZoTwJCNLL;\\\"\\\",2):f(\\\"\\\"{bn5B25zhbbuYG,l\\\"\\\",2):f(\\\"\\\"{qSBE8<aTaFa4pFL44m<ujix-\\\"\\\",2):f(\\\"\\\"}AL7rFL2q<zuCTaJC4.Fi>,Hyx3K.1-?6?-h>d1>6O=8,YaB2G2C-WZ;+P|izGij|WZI5:AJ-n5jbA/DagbhI2b\\\"\\\",2):f(\\\"\\\"{HSin5UwFqGI5HpYN2J-/bEaWZkb6b@tHy=uLV/1s3agaNDYa7gr4/ea.b?<x6exdFaZ03bAf:z+:3<Oz1P@a01588sYYfO+bD84b<,EDG.\\\"\\\",2):f(\\\"\\\"}b;pgpmO3zopXay5y\\\"\\\",2):f(\\\"\\\"{:3GES28zopkMZuJ<S/p<DalJjbxUw\\\"\\\",2):f(\\\"\\\"}tb=uTy.>RGTaibdv6WDaXay5sTE7I*Tr*8wbGhQIv*ubkb=QOaY*Uvgb8buj6YfbebEcxpfM:u2bWalJDyc*hb8|pO;RCzxb5T3r01j,GN:zv|i-GPEavbDCbPiW=z-Hoq75Jw<ag"));
$write("%s",(";gbFaUv9Vp<W/CR|bH\\\"\\\",2):f(\\\"\\\"{zpjb|K\\\"\\\",2):f(\\\"\\\"}bTUWaIhtbpOrQcXBr2;35nIUq-dP|B\\\"\\\",2):f(\\\"\\\"}$6ezdXay5wbD@A=1p7bOt|bYEVSSoebabE0sx,3+b3bwbK3RDa+0Albmr9;3:W/CRnXkb\\\"\\\",2):f(\\\"\\\"{bMh|BM?nSRtS\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{dHUIh|bdbMY8\\\"\\\",2):f(\\\"\\\"{8b+t.bUAJ,aBiu*VB2ENub2+/r-TwxbUL\\\"\\\",2):f(\\\"\\\"}cj9wp0:x01wb*bfbNazpCaNaw\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}9d5FhmsFatbQ0mMiubb8\\\"\\\",2):f(\\\"\\\"}oL4\\\"\\\",2):f(\\\"\\\"}wH*BDaUCj\\\"\\\",2):f(\\\"\\\"{S4EG\\\"\\\",2):f(\\\"\\\"}Yv9Mq7K4s|pUv3gSRDBabAiK4N2yEA\\\"\\\",2):f(\\\"\\\"{BaewtbybkbK41ba7u6dbK>\\\"\\\",2):f(\\\"\\\"{>\\\"\\\",2):f(\\\"\\\"{u1bJ4eQ\\\"\\\",2):f(\\\"\\\"{bRaj*>aL3Jq\\\"\\\",2):f(\\\"\\\"}HUCj\\\"\\\",2):f(\\\"\\\"{?2q5rI:\\\"\\\",2):f(\\\"\\\"{D>lA&6e.dAahbGafOjbsR\\\"\\\",2):f(\\\"\\\"{DAYxB+5?auFK3/wO?0b7bSc>aKoW/hQrDRuPw1\\\"\\\",2):f(\\\"\\\"{dbiiH1/b=,\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"fbb\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"}LV+bwbebzbHHPa-bS/9wvbK<yb<aG,k=x24U;,sCh0m*RWebYYL=C*qskbOXp+>Lq*NaG8-biiS3vbBr2x>a<a/+p\\\"\\\",2):f(\\\"\\\"}zbX*w:-xED<ax,XxZ4/b<,l+dbYYbY<,cCN99+|I8qDCE\\\"\\\",2):f(\\\"\\\"}wbRG0|N|t>FE>ok<LukbTaNDRaFatboNwb:,i/f+6S9GtJk;2zqs8>Va8bDaejs9ej8b2b0B/r70vb;tUZiilVB2j-88\\\"\\\",2):f(\\\"\\\"{Gtb@aa-oOhxdInSybPa\\\"\\\",2):f(\\\"\\\"{bTaB6Pa22-HoqP<3ugu4bKo>afbr*trDa\\\"\\\",2):f(\\\"\\\"}b:PB4Um6+3bQv4JGxVxLSgOb3OF1brU,b1ba>kzSZs;\\\"\\\",2):f(\\\"\\\"{qj,>oks?af4sHh@LuI/*bxsN,W@H,l2p\\\"\\\",2):f(\\\"\\\"}nxRtwHgt6b?S?-0:tb6>UaZtVttbxhii=<Q.+bDBtvDSeb|*I;GyXa=.;voXt59TUDv.sHYh>Yub4yqr4pZrsEx+6btULzj/OaG*uw*|X8zbqCI,KrS32bWa5qs\\\"\\\",2):f(\\\"\\\"}<X:\\\"\\\",2):f(\\\"\\\"{=stG0ANaM7Eaibgt6bIkdburI|XzUrkr58l2wfDfUaP>,pRa1bn6:JUrYo22FFUr8bujUttb7x24>.\\\"\\\",2):f(\\\"\\\"}z+t3uUrRIqQW?UqWaGRVzlR=Qlb;,\\\"\\\",2):f(\\\"\\\"{duwE4R"));
$write("%s",("=V9RtABd6a9aA*9zBqUv\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}v1P\\\"\\\",2):f(\\\"\\\"{qC14kbgsjb-bW|i\\\"\\\",2):f(\\\"\\\"}zptR|bii?NFy;j?fG8DHVad4a<bGF.Be3zMQ?\\\"\\\",2):f(\\\"\\\"{3t->|c.8Ct-16GIgbgb>aP\\\"\\\",2):f(\\\"\\\"}/u0:hbxb3Lf9=re\\\"\\\",2):f(\\\"\\\"{e9.bnXkb-\\\"\\\",2):f(\\\"\\\"{0:5bNa4sqOv>u-7M+3rgQwFw\\\"\\\",2):f(\\\"\\\"}bn3a@iFMv.b=r/uLQiiyr\\\"\\\",2):f(\\\"\\\"}b*b=BX.2bUqIt?6\\\"\\\",2):f(\\\"\\\"}bYaf0S\\\"\\\",2):f(\\\"\\\"{fbgbRaa:OS<a-UfBg\\\"\\\",2):f(\\\"\\\"{+dLt0;XG5I24=0NaX.;zfh+rWaDav/DaYhuFrDPiEM.bQ5N,\\\"\\\",2):f(\\\"\\\"}b8tPa2bz?:>-TjEabT;k4?6QafM3b\\\"\\\",2):f(\\\"\\\"{B=uldwb@uPvfbEaGafONuE\\\"\\\",2):f(\\\"\\\"{p|>\\\"\\\",2):f(\\\"\\\"}vbab0BO8.bh+P2WZPa-bt1:,Z7;p7babH2TaDqjX8z4pq.SY>a@ucIPaUa=qmyG6E68s4wCrbbz\\\"\\\",2):f(\\\"\\\"{x\\\"\\\",2):f(\\\"\\\"{|fVavbPr2bn*uFK3?6PJ/*|tp-@STa5Jor2t@tRoNT5bZzTan0mJG,+0OXo-nMz-QuCrPa--i/2b7w+-w7|5f92p\\\"\\\",2):f("));
$write("%s",("\\\"\\\"{bTaFa.bZa?ap;as5s;M-C0G0S\\\"\\\",2):f(\\\"\\\"}yA0*|Aa=au0/@>au*mdk|S>Q.r\\\"\\\",2):f(\\\"\\\"{Sa\\\"\\\",2):f(\\\"\\\"{,@.c.w\\\"\\\",2):f(\\\"\\\"}l\\\"\\\",2):f(\\\"\\\"{J2u;4\\\"\\\",2):f(\\\"\\\"{No:>|sOv,2u<6qbbW5wbpDnD\\\"\\\",2):f(\\\"\\\"{blDUaJ*Y7n3Qi-TnMu;s<t,X>hb7bab/bCzTa4wmQRa;A@|EqFTaL*--nI\\\"\\\",2):f(\\\"\\\"}97Ko15bbftx:SvM<1\\\"\\\",2):f(\\\"\\\"}RBu<Iqvb|DJCFGiistkwRDO=O9ybcCn,sWrQBwFDss29Srn,?t;v9vOWk|n,hujb8bktE:*Va\\\"\\\",2):f(\\\"\\\"{fs/uLQKfkboNEaPDlbVQabc*tb/AD@7brq+VTq+5Ga9W+Wv>@aYaMvk2Dqx5OzK9e|azp=0UxJDdUJDXx=0Y;Tas3Q?:o0sEf8aQaO;d*<a1\\\"\\\",2):f(\\\"\\\"}HUf0E5Z9PaybZ9UW?GtbwGp\\\"\\\",2):f(\\\"\\\"}hbtb>aM,-xCyhJ?iuhHb&b*2x<nI9w6b5|n+uw6s8ZgbgGcDebB2=a;qLL+0@uZC0q:A*bk,Gxm\\\"\\\",2):f(\\\"\\\"}qQm9l\\\"\\\",2):f(\\\"\\\"{-.i.8AOA>awb6p?a1bL+kuKxh4EaUT4iALXWOu>|>acy\\\"\\\",2):f(\\\"\\\"}b,:|by@|/:AZBwbw3cAaCI013ujqZCP\\\"\\\",2):f(\\\""));
$write("%s",("\\\"}s:gx;-Dqfm,:LV|.o8G,zdJ-m7,+B/TC8H0sjdWAldy.*b54$6eHbhHNadp5>p-4opTib\\\"\\\",2):f(\\\"\\\"{b1LF-|ya/<aB6-b|yU-:um\\\"\\\",2):f(\\\"\\\"}s7VaRt1tN,I:*2UrUqm\\\"\\\",2):f(\\\"\\\"{ev.:d+QJ/=aVkbW4FavrybRac*l2PaOa:\\\"\\\",2):f(\\\"\\\"}?aE1Da5.*sqCE4q:QTUv,4<aybIuYar8nt|Bds9wk4iwp+7bPVjwFaDqiiH1+3c*b,s,|ybZQd3hVK?oN=;*b8T?iO;jWqrzpIqFavus<1s;slsNxrV>WRa-A+bN9A8p\\\"\\\",2):f(\\\"\\\"{4U;;CRPJ.w/rX4vGA\\\"\\\",2):f(\\\"\\\"{jb0b|w?GswtbX0a+du2bkb48tbirQoqw>a/waUguBq&6eqa5.EXqr78-A@|ktBqo3a2b|w>aRWujd83rKU0=Pa\\\"\\\",2):f(\\\"\\\"{bC\\\"\\\",2):f(\\\"\\\"{01\\\"\\\",2):f(\\\"\\\"}bN*ylUk/|U3AsC7Wa@3=5:2EFnLUai1?aA8|QN5aOiu+pWNm=San5zb*.\\\"\\\",2):f(\\\"\\\"{86b1BuF9ba1K4;Bm<?qBpd*Bpv-g59Tn3Oa\\\"\\\",2):f(\\\"\\\"{bjrn5z6Pao81bi3aCag:tv@adsd5|z5q<a<aOa7btR.b8bgvfbw\\\"\\\",2):f(\\\"\\\"}cb5wy|mpN9hHvsYEftNx|HZa@axri3ama6bD2UanUPayX[3c^1^\\\"\\\",4):f("));
$write("%s",("\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'aVaXatv@aax7bn<H..jp*=z6sI,1b*5xrKU?Eaeajbtw8@e|b/w2b/bkb6\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{79bCrfbtBE:hb1bBwxbBaE5K4v-tREa7B?6RakbXW;;X4RaJdybnIQi?2>|GjbbybX*a1dwrxBfQ=\\\"\\\",2):f(\\\"\\\"{b.vZ?xvi*RBccoSK/RWzb.vvf\\\"\\\",2):f(\\\"\\\"{KaWbDqDBCkEUcbRL2v*BwhOYK>JvwbYFM|9bxbibCVzTdbub+b6J4p<aRWGjZa4Ijb.wVi1r<aX2ldOu6b\\\"\\\",2):f(\\\"\\\"{b:xcvgN\\\"\\\",2):f(\\\"\\\"}w@a;;:,/rX4R9FSjbq2zbgp4w@oNa\\\"\\\",2):f(\\\"\\\"{bubcbW=k,w.Er?ag;;LxwvsIuvsDN2vE:rIj\\\"\\\",2):f(\\\"\\\"{vbrqR0,bGa>DvbrS9fxdR0/xL,Na;+2bKU?mlwmbB-l\\\"\\\",2):f(\\\"\\\"{ab*-.0=udxAukzXaL<3b:u8u\\\"\\\",2):f(\\\"\\\"{dr1=tPV6=Ca+bybdbfyGKqw"));
$write("%s",("f;4B+p,z=uzS+x6bUk<l+b-ur1*?|/A5G-ZrdSHJs;L;28@u6PIy>a/bkbC;A;<s0/pqRz2=gb8+o34ikbjvebXa:\\\"\\\",2):f(\\\"\\\"}-zQaoD0skrUDPvFavZP|hb;tE0sxfc?Gmb6P0@cI6W/=3b\\\"\\\",2):f(\\\"\\\"{<xbYa,@c.O4d.UarM.bAuaV:Arxt3DyhbgpRQZpWaGjxxIEb.Q.DI:8DI?<iiyr2+p-5b>8wbIC$6ejb9r8ZFa/ub@RaX2vb7qEaiiQJfb@YyQGafOGx+38b-b*r7b0:\\\"\\\",2):f(\\\"\\\"{bOwRu9AqKBaix78Q.0\\\"\\\",2):f(\\\"\\\"{-d9x0:\\\"\\\",2):f(\\\"\\\"{b5bffmbSUeQOa\\\"\\\",2):f(\\\"\\\"{b/^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fla\\\"\\\",2):f(\\\"\\\"})36(f\\\"\\\",2):f(\\\"\\\"{#,43z3m|a7693(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})8402(f\\\"\\\",2):f(\\\"\\\"{#)K34BauB|Qa?<:o/HEQ:jXW>0O68bhuk+N\\\"\\\",2):f(\\\"\\\"{iHt@/O1bYap=ATk1DqO6XYRrpsx2vwaLpYe-bjbQaGsrUAiVKU7wbiUK5/wH5<*Uv+QvM,=G50g@av/6@Y5dzLrVaI/0g@alb@@>@n\\\"\\\",2):f(\\\"\\\""));
$write("%s",("}U?MM>ai/\\\"\\\",2):f(\\\"\\\"{bOSX0LMQ.DIAsSOe3q.ow8bi5ibCaX5tPm=b1e63PPrab0g@pqKSHOfbblbUtt1>atbzcYaRGlbOSJ@8be3>aN.bc5-Va0<6rS-YS?aN\\\"\\\",2):f(\\\"\\\"{i5r.tb<,;B?vEa;3mbv2*uIQt*Dq27lbUtV8qKR-o5a\\\"\\\",2):f(\\\"\\\"{cRaW<Sa<jB|YBsFe3G5ZaGicbiq*vvbXrJ2S4\\\"\\\",2):f(\\\"\\\"}HM.GxrD1Xubf?z*Va8bUvB4UmXo22|b*BkbR/2ze\\\"\\\",2):f(\\\"\\\"{Taa@nLfg\\\"\\\",2):f(\\\"\\\"{HzwSATWRaF,Na\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}nEUaRa1bX*iih44LO.v+Rtfg8HN\\\"\\\",2):f(\\\"\\\"{oO@zm9*CFT;t-v15Nag:Uaj8t1GaFT5bmbN515Na90BaR9fb1bX2w3kb5b7bF72K\\\"\\\",2):f(\\\"\\\"}qS4\\\"\\\",2):f(\\\"\\\"}H.6e)c6PXYibc\\\"\\\",2):f(\\\"\\\"{cvmyIGs\\\"\\\",2):f(\\\"\\\"},l<aKuXaBzjbRLmbSUgretOWb@.b4z*.>a8bG@8bDaiiS./b6>vbPA/|GjxxjlY7g-+xc.u6mbpXdb\\\"\\\",2):f(\\\"\\\"{VxXFMZ:cbJ,|t<oSay.4oDM-2Q-Nay@vv2vPa/bQ@6bRaWhtb\\\"\\\",2):f(\\\"\\\"{w1pVarDebBR6q77K>o3uLQa\\\"\\\",2):f(\\\"\\\"}-nRW/Aa"));
$write("%s",("QaPajb|tI/NaiWU-P<JJg8>a0hbpbvhp4>|4aQaRaySa.Dqkb2qOUiiQJdsn/Xrr8-:eb45OwjXG/.2b2lNRzKt9TlpiF;;*2\\\"\\\",2):f(\\\"\\\"}bTaRDTwb@BahMi.Du,6e+a\\\"\\\",2):f(\\\"\\\"{b.QP,l5w\\\"\\\",2):f(\\\"\\\"}5bhbPR7x1b7bU3ZaVx/zk2Da6:N\\\"\\\",2):f(\\\"\\\"{D4aBc.bBw1ia1*bVv-4C.nSDqN5h2l|A-u|WaKUU6gbUawsUaP:ztldqAz3228+Nr.bnv40KtsYab\\\"\\\",2):f(\\\"\\\"}*Z\\\"\\\",2):f(\\\"\\\"{2bY7*dZQ\\\"\\\",2):f(\\\"\\\"{DdbZa8qv<*.Q<ib+3l:R6wbCRjFf4X|.,x/1b|bS*EqbYnIE:@\\\"\\\",2):f(\\\"\\\"{8XdwCylb8z78tvx2kbQ=@aYak,ztE1,lj|IMnPax>,vGAajva1t0MIh<3jZa3trGguoFZadbAs,sm*qQW?V5WaI6RD0=bq\\\"\\\",2):f(\\\"\\\"}YUq64Ef|bTLs|v9dwZaGu?;R=sY+?Ta\\\"\\\",2):f(\\\"\\\"{DdbjnvsFo@qldBr9;*5UkmP2IBa=a2brx\\\"\\\",2):f(\\\"\\\"}CE9Za3rp*wx<a=aV|Uwmutvsw58fpubPRhJPa*bNt|zk4dbALtvCN*b.|?3csa77Sav9E9E:Io\\\"\\\",2):f(\\\"\\\"}CIgQ=\\\"\\\",2):f(\\\"\\\"}Ha2b*w6bfs22Ta-.xhqRTw-L-u*LfwL,3tm@\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"}6xbUCWaz6Tajbgtet,3z*z,Fi2IlJRat0t|ftX>|t?mlCRIlJ>ads?-Z0iCe,|>?mFai\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{36NO/1BaSZE7Dq=.guOWSRU68Hcyz6e%dA-OWDIhbnRFabbDq?s3bt-djSrVaj*>aIHyjpGS>c9JqDqO?TaibHrhH=albCu\\\"\\\",2):f(\\\"\\\"}bKFSxtxqpMwc9|bcj2pW0uRs9\\\"\\\",2):f(\\\"\\\"}b|DEnt0MI7qmhh<3jdb>322TaI,\\\"\\\",2):f(\\\"\\\"}:FVnRFaTrA3cb>jAa-bt1ybWt9A7-hvEoGpv2?aVtX0p<lbLoHRZxL\\\"\\\",2):f(\\\"\\\"}jbQa<.BrufLowGX7|bkb>alxzSiC<a3bMRixD1v9lIbbEUH\\\"\\\",2):f(\\\"\\\"{TBbb-rvFScBas<-bD31lyw<awbXaCt0;\\\"\\\",2):f(\\\"\\\"}Hcx>|zBp;N9\\\"\\\",2):f(\\\"\\\"{uN9?8AaNt4B.b=.Va@p4BpXj.CuChDfbbvFxb*uHraby.RQ9r4By.Uq/hBa-sSaoq>2Sacz6o@q4B/h8.Bac\\\"\\\",2):f(\\\"\\\"{+b0|.d7M8.n58.8ZzbSawr2s0|zbvF.dXh9;;3a[a7bzbUa>|oTcbPRlbGabY;sCzpSCzGRSaEn6=hDzt-N5|Sa>P<Zp:<Zp:ybyJwb*.p:ybIx\\\"\\\",2):f(\\\"\\\"}b*.p:<ZtbeVzCFFc3apbO,P5u\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"}Aa>aP,yb58|shOyJDqGpgbDLEa-bzS:\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{85bnx;3fhHsYzVt1:,sL\\\"\\\",2):f(\\\"\\\"}Iq\\\"\\\",2):f(\\\"\\\"{b4ibbw\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}w5bqS-t;;v>TaIqxbyuJzyuu/PK+sA>(6ezcesauIQqregirs,@SB0wuNa+1w\\\"\\\",2):f(\\\"\\\"}/wjX@6eG-W@zOwUa=+k6A3?p,si\\\"\\\",2):f(\\\"\\\"}6bPaTBZa@9SaibHRfIS\\\"\\\",2):f(\\\"\\\"}iUo1L<n*ev5bNaL<.bkYCyqS-tLGNa;32be0UCfyv\\\"\\\",2):f(\\\"\\\"}wUp*?q45r>XaPUlsP3>afb;rG<Q<6p<agbR|W0;3fgbThb/w\\\"\\\",2):f(\\\"\\\"}b0;tbmPJ3-tGr.b8,fbUaI652\\\"\\\",2):f(\\\"\\\"{D5w0=>.0/KdSa\\\"\\\",2):f(\\\"\\\"{>\\\"\\\",2):f(\\\"\\\"{uKfDaeQebRWC<E114t|jbdNT2htKj>aE114Gi*b?@xbr17zv1F;WacxWa1p1b2b/b=uWaaqr8oK&6e,b|b@r-NBa<acbE9y\\\"\\\",2):f(\\\"\\\"{n0|z@iw<T-s\\\"\\\",2):f(\\\"\\\"}rx0*;\\\"\\\",2):f(\\\"\\\"}yw/+AU3LX0RCEPZa@upM>wn0W/k\\\"\\\",2):f(\\\"\\\"}N.RaSZEDPa5b4\\\"\\\",2):f(\\\"\\\"{?qhbv9TaqzOWy@a\\\"\\\",2):f(\\\"\\\"{-"));
$write("%s",("bR\\\"\\\",2):f(\\\"\\\"{<a5.E:*|\\\"\\\",2):f(\\\"\\\"}br1|MN+cw7b*V7-PvRA?aD4aBbk8RIqQ>07tgbXa<*Uvv/680@>q-bT2gv*.6@RoZa7gn|Ca\\\"\\\",2):f(\\\"\\\"{bT2uqOF/xbRBwtK\\\"\\\",2):f(\\\"\\\"}bpsI:XXbbibRGD@/|f\\\"\\\",2):f(\\\"\\\"}8L+uL<fyjtJnPC=o@pUmybUH?21bgtetUmB\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{|bGA2b,|g3RavqvbZa64FuN+E2|6ehbnweQ7b>SC-nMY5gb89LNoXR,DCO,z>6zSOP\\\"\\\",2):f(\\\"\\\"}@a.b7tF+7bK5VaO?i-Q<k2W2V8HdGjkbGhjbB?WoXYu9zpw3kb2ICWS.o4K7a>blB>Wn|FzOq;,Lhe5Q4Fa0=?GDq=aTajbPV/klT8bb@.bj6H>gIqKv\\\"\\\",2):f(\\\"\\\"{UWgff,mbNuqz2zuuu<dbsYq>sz>?r\\\"\\\",2):f(\\\"\\\"{8ZIQM/wt\\\"\\\",2):f(\\\"\\\"{bOw?:?6>NLjgTtviUGXkT@uE7ey88@qZa*b<,fbfEtbE77b\\\"\\\",2):f(\\\"\\\"}790+3ara525|I,;A\\\"\\\",2):f(\\\"\\\"{*Du.j?6E)3da=fY2yNyC-iws9fbVJubeb:2=x40Ya:t8tGaV3wshHSa0sEa5L8bbU,u\\\"\\\",2):f(\\\"\\\"{4DZkY90LG|F4b4Mi37Lm<90EN\\\"\\\",2):f(\\\"\\\""));
$write("%s",("{bcr5b40fbjPFavMebPvRWwbW*449by>;t2U.d>sl>FG,tJ4C<k\\\"\\\",2):f(\\\"\\\"}Q.=Bf71;6qdw\\\"\\\",2):f(\\\"\\\"},IC@qB\\\"\\\",2):f(\\\"\\\"{kR77/wN/C.msZ4C,=Y<axbF;p+GaEYoHj\\\"\\\",2):f(\\\"\\\"}FLlWtbF;y.GaBWq*dbjKhba1SB9sjDiiupN9n\\\"\\\",2):f(\\\"\\\"{kYFafb5LT+q2S/+:nt;wxs9slb6q>\\\"\\\",2):f(\\\"\\\"}j>wxUqjbdzu/AB/bpYEPTah0|Qa-1SxW.GvWyy*W\\\"\\\",2):f(\\\"\\\"}b9;:okYn0jD,bOqYaT\\\"\\\",2):f(\\\"\\\"}Qw.B.,,lA-a5iirL=ag;I,CO2GUD+bR9F,9pKq\\\"\\\",2):f(\\\"\\\"},*bIwjwgcx22gv;pwBaY7Va@*lA+pn,;F3xdrZavbwqnDf+|bq8n5ICOrQDNw,z/wTrmbybXs;tbykbQcm<-NVa=aFaHS-AqshuvvtCSa4b4b\\\"\\\",2):f(\\\"\\\"{=\\\"\\\",2):f(\\\"\\\"{u\\\"\\\",2):f(\\\"\\\"}bSa?<g0vbB8<a?4-b<a\\\"\\\",2):f(\\\"\\\"}b,bQaybRSPaQaXaI>7bu61L@a+1WadNPq8b|rBKj|\\\"\\\",2):f(\\\"\\\"{u\\\"\\\",2):f(\\\"\\\"}80tiiTvLj6WLS<a4icj1iu@MKdwGaD=ls5pS4+vOavs@vwbFaxn3bbb4TA3FOyi>ML8|A\\\"\\\",2):f(\\\"\\\"{UabeVXaY:mw8b/+Cs>Ub"));
$write("%s",("bguGu6bDq2gl5>ygp\\\"\\\",2):f(\\\"\\\"},IUI,kbRappQzuV-,hDT4fmeb0bqLY?qz7bjr|OUC|Ny9ybGq4b=a1by:YpnIED5pYxCrF,/r/09JHqt1e@Tw/|U-xw0tBss<pQ-x+bMI-A.bxb.r=TQz*bcx2-2babw:RaOz9t7t*L?Gwj>3XaE5Jwdb0soN5|ubyEWU7\\\"\\\",2):f(\\\"\\\"{SOUqmbebG-zw1ptb2bb+7r?G5bM/vb7bSz<r@aC<ibkuE:Ipii;5?2Z\\\"\\\",2):f(\\\"\\\"}2q\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}UaUTWhGac++bV+hb\\\"\\\",2):f(\\\"\\\"}@9rqLDqSr>Rfk=K0CK8/Sv,Nyp*dUt/6sXaixdbTOGFL5c/Hqp0rGvrgbaPd5uyab7bZt1bhbsRqsE\\\"\\\",2):f(\\\"\\\"{Urv,cbMQQazbRaybZ\\\"\\\",2):f(\\\"\\\"}3b,+eTy3fS.7IdiirTh2lws22D;,|<s2Xy|btuCNPtwbTanE-p8A<a\\\"\\\",2):f(\\\"\\\"{dQS2;y,b+x5Ba\\\"\\\",2):f(\\\"\\\"{b@a/<7oWJ.j8brxgDQ7Qwm2ebt>QaX<Ra@a,</t?ahHR\\\"\\\",2):f(\\\"\\\"{u9nQPahtjb/2vKDSO9nEJ5CcMIdbiuU6@aib|bKywbcba>ubmxj6D\\\"\\\",2):f(\\\"\\\"}vbHsnrb+7bARvL:Sxb\\\"\\\",2):f(\\\"\\\"}9*beznHv\\\"\\\",2):f(\\\"\\\"}o|5gYacu3by+gq"));
$write("%s",("cN-y*A=M2Q1P2\\\"\\\",2):f(\\\"\\\"{Ratx<*b+DaNawbDqWvjnSOUar8Mon/0b>aub\\\"\\\",2):f(\\\"\\\"{bq2?p,tAag8qC-9>aRA9JlAqLabQ@Lf-/f\\\"\\\",2):f(\\\"\\\"}qLQ<kuDqW0N+tbp\\\"\\\",2):f(\\\"\\\"{fb0qe5H|+by+0b,b/|9bCs6QNab+kroD\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"},+xL>aX6I6t|z>cN5uiCjv9syu,bgGJ-pl,2z1uwplPBW@kKRzP0Qir*hbubYaI>ubmvY*Vat:?afbfbkriw\\\"\\\",2):f(\\\"\\\"}b-bp<P0i*JoybTaGo9rqQXE9zXaGuwbB/4b:Q/u3b\\\"\\\",2):f(\\\"\\\"{r9bO=|b1KeG\\\"\\\",2):f(\\\"\\\"{?9bR\\\"\\\",2):f(\\\"\\\"{i/aq.6bbqADCxbDw?q.bhbzbiiMtI>Oq;M;O6+9z4ps2;zfsv2vqQ0qpard11\\\"\\\",2):f(\\\"\\\"}Hgbb*,jtSIYztbfb|bn<EaML=Htu:rGaXI8qGsVaOoQrcbk\\\"\\\",2):f(\\\"\\\"}+bUH4q2q0qWqkrU\\\"\\\",2):f(\\\"\\\"}tAroA0j3SG<7vq?i=r0;=zm/fsi<6px52i5b9blsfb|pDa|4t>:\\\"\\\",2):f(\\\"\\\"}B\\\"\\\",2):f(\\\"\\\"},@tb4HxbEaKhTa6pI:Kw4w\\\"\\\",2):f(\\\"\\\"{?K\\\"\\\",2):f(\\\"\\\"}4e5+C923tplp=NSr,u4/Wamz?=:D/ba:wbdbX>5b|"));
$write("%s",("bG9Ba7bvKT\\\"\\\",2):f(\\\"\\\"}whQ<Oa6=@|0NE2-bYoIBLM8blsp|n|?elb;qy9UC;ux+HhfbWIc\\\"\\\",2):f(\\\"\\\"{roFaK\\\"\\\",2):f(\\\"\\\"}Ea-y>//Gbk.C;MG>;u<+:+my9Mt05t8bxDUaCaTC4b<a+LmClb6bybAaE2Fahh/bTwq>a:W0yb.bdbF;Aa9b-bO-E:QaiiY3>ycN>+?abb|bb6O,h3Qa4,Q7LpDaf8-u4A\\\"\\\",2):f(\\\"\\\"}bP,+b\\\"\\\",2):f(\\\"\\\"}bXa2DFFUa:uybjbSaE\\\"\\\",2):f(\\\"\\\"{90c36b:NGq?6pl8zhb\\\"\\\",2):f(\\\"\\\"}bOw*sUoZaHr01DKdb3bfv\\\"\\\",2):f(\\\"\\\"}bmbj,\\\"\\\",2):f(\\\"\\\"{092-bUaXa|u>x-,*F=aDK6xabhbBs\\\"\\\",2):f(\\\"\\\"{beti<CaCu8>s<k-XuH>>+ubUaLGQ-B=e*ZuWa8bk|DIJIS>XkS>e6p,;uUaB<-sBadsN<MLWaSa6rF,*7yyiks?<K.y:Keb\\\"\\\",2):f(\\\"\\\"}4;;fbtb?28b@vRtH5i*9Hl,/67q2iUJ\\\"\\\",2):f(\\\"\\\"{,hb8s:3tKF2xD<a+bUv@|;tH\\\"\\\",2):f(\\\"\\\"}c:y78b<a@aDq<a7.FaFjXaXEKtr,XavbQaN5+55-+bFaOao|2b7bf9H5@aUa>al=j=z?D8>aDaG6kb@@N4Daf\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}qkb3zfy8;58i3"));
$write("%s",("ZaLv0bq>?a.bUm|by5UxD3XC5bFg/bt-|016Ta09xbE4>aQa?un63bPaXa6\\\"\\\",2):f(\\\"\\\"}Ean5B/bbM?Qa?s\\\"\\\",2):f(\\\"\\\"}636hzI>y+tbAa>rfvi\\\"\\\",2):f(\\\"\\\"{R\\\"\\\",2):f(\\\"\\\"}UaJoiz=a*2Lo6=\\\"\\\",2):f(\\\"\\\"{w<58bEHebGjXrHrVaDq+7Bau/s,=mx\\\"\\\",2):f(\\\"\\\"}?<S1f=:I</5E2b;\\\"\\\",2):f(\\\"\\\"}IuA3hpV5L<,b0:kEDoEawADqk4a>GaY=RaW\\\"\\\",2):f(\\\"\\\"}Bah?db1bKuUk:|gbQal@,b-bbH\\\"\\\",2):f(\\\"\\\"{IFuVakb;tgx8HB2Gxqtr6u>Nxo>|58b5b?aduoivs.b0bUA4bHIR,l/tbS68bn;euN/Dc=sarqJlrIg=.u9RImxm7,bQqTa7u@a\\\"\\\",2):f(\\\"\\\"{bj/4bo4M>5;Sc5;2bybIBFaCa=qhv<aH\\\"\\\",2):f(\\\"\\\"{/=DIM<rgpp*bcbhc.rIr.bXax64+WA?a?qSvlr.-8b88.IFaiiU0Ya=.fbSaybVa6bMv;@>-=ae3P>Wa16/bWaAzR-QaVaK4J9eu\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"ubK-=s-y1C7IS:u4+GddDahbT6Ea>3619bSa+d.qY;S-yyA0i>c;r.?pwbkArxUCX-ub5boi\\\"\\\",2):f(\\\"\\\"{bjbbli\\\"\\\",2):f(\\\"\\\"}@\\\"\\\",2):f(\\\"\\\"{WF2z:uebDqXv44x"));
$write("%s",("bWw5,oim9RaRGGa0HJqc?u=rqE\\\"\\\",2):f(\\\"\\\"{tuS4CaRG5bFaRa?au\\\"\\\",2):f(\\\"\\\"{TyUap<\\\"\\\",2):f(\\\"\\\"}b>a/Hmb=sn*>aa/Pzy\\\"\\\",2):f(\\\"\\\"}QwZalrxbb@lb=smuiio0<a7bPa.q4ocbzbmbJ-;@E5=aiba.2G9Gu<DqRa+bLofbRa<lF*AaGa:Fu6bcvbnt\\\"\\\",2):f(\\\"\\\"{.c?v2X7*bQa8q2sX*Cawb@aFgyb.+M>V\\\"\\\",2):f(\\\"\\\"{ebkbftBaZC=ayb?ajDt+rD8Gi\\\"\\\",2):f(\\\"\\\"}FaSaxbjw2b60zbybAB?p-nE:<a/bfk:/\\\"\\\",2):f(\\\"\\\"}AS1\\\"\\\",2):f(\\\"\\\"{AV1yAU,n*A1.bzb>a>,RaC6k;-bn0db5|Va>pg*k4Cy+iotDyMqbbCyzbc\\\"\\\",2):f(\\\"\\\"{,rNv6bE3a@=a6pFoab2wZaUrAso|,bIpNxhbTa5,HClt4bdbzb854iE53bWaebPaA5eyiifz<|,qyw+bWhI5\\\"\\\",2):f(\\\"\\\"{Bz/896949D>u9Bfh;f;ov\\\"\\\",2):f(\\\"\\\"}b.D6b5pe?s-D3bbctWa-xv/hblbY\\\"\\\",2):f(\\\"\\\"}ur*?LtJt/b4y>+OuQ.Ihn3m<kEU8eb+b|fqAfpJdiilE,bz*5b2b;+@;9=krVaqsGxPa9bV5wEq:Wat,K4h?jzP:Ea/9F6cb8ubk3ETn,C,4|bvbb@n|I0-:4yr1b?B/\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}67sTaOvMC154s>+Ca0b=ouBRaPassbbFa\\\"\\\",2):f(\\\"\\\"}b82pxCuWaix+9\\\"\\\",2):f(\\\"\\\"}9j,K3FazbPcB|0:abfbbb5b.b\\\"\\\",2):f(\\\"\\\"}bjyXaubbvTaXaSxj*hxOaxb*bbbIpY\\\"\\\",2):f(\\\"\\\"}exiirs\\\"\\\",2):f(\\\"\\\"{b0swwN*8b;?E0n56j09Ua,b+qovLvBxP=Q94C|DQ-1bUaDa@\\\"\\\",2):f(\\\"\\\"}mbv\\\"\\\",2):f(\\\"\\\"{Nt/qv7HxTa\\\"\\\",2):f(\\\"\\\"}4W5cbmb,*fbv7TaFxibFap,*4Qa=ab.iq6bO?<a=uzd>acbW0Qau,4bV5QzczP5:u|b/b,+kb36J3Fa,2ib6|ZAsBhb=aUaZajd.s\\\"\\\",2):f(\\\"\\\"}bi/70lA,b/bVp<6t4Ssp?ikn?vyGa03-x\\\"\\\",2):f(\\\"\\\"{b0bF8z25,<t=a.bX*8,Za63Q\\\"\\\",2):f(\\\"\\\"}5s*bH\\\"\\\",2):f(\\\"\\\"{2b\\\"\\\",2):f(\\\"\\\"}++bO\\\"\\\",2):f(\\\"\\\"{Yx/AFaWA5blwMz\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"}b/=J3Q/F,Va<aNaAaybDqX0C<lbpuLA9b+pkbi>QxOag+fhWaYa/bv+cbh-5bDa9bzds2fpm\\\"\\\",2):f(\\\"\\\"}abF22bPa.b*,gbVa27/s/bC7\\\"\\\",2):f(\\\"\\\"{bhb|bXvLpJwJ*Da79q>mug+5b+b\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"}\\\"\\\",2):f(\\\"\\\"}d8,bdBqrC-?aNa7,/w8sx+g;W*5bUm.wNau\\\"\\\",2):f(\\\"\\\"{kboAebibDaCaVa|b2hYy40E:c8f\\\"\\\",2):f(\\\"\\\"{d\\\"\\\",2):f(\\\"\\\"{,bp*:>1\\\"\\\",2):f(\\\"\\\"}ebw0uuSvK9vuq>Aa0bbbYa5yUmId-b?r25Y2\\\"\\\",2):f(\\\"\\\"{b6bvblAXaRtVp5*r?a-J8Cvw4/dQabcewPzPitbXaguNaDqXa-bBaP>zr|bYa1tB65>Wa-bubM:u=54Oa<aWaE3z,4\\\"\\\",2):f(\\\"\\\"{8bl,wxXaGp-qi5k;i<hbEa77D|bbn@rp<@EaRaf;;3Vt@a9z:0dsv2mbX/i5:.x6-b*bVa9z\\\"\\\",2):f(\\\"\\\"{.Oav/1iq>D1u\\\"\\\",2):f(\\\"\\\"}=ambO,wbZ9ii6mhb;8J2p-35xbCa=a3bbv90kba@\\\"\\\",2):f(\\\"\\\"}ugbgcr6gb5bSaRai<5bPoxbu\\\"\\\",2):f(\\\"\\\"}xxOaCaSa|b8b8b6>4>Iw@352\\\"\\\",2):f(\\\"\\\"{?52Eaj|8odbsux;3b7bGx07Z\\\"\\\",2):f(\\\"\\\"{Bovqn|6bI3Sa6y:\\\"\\\",2):f(\\\"\\\"}3j|b28Bzld4bc*,bhb0wEambtb/6|>lb:tb6fkg|e=ikc=fka=bbN5qrZ0Zp?u55xwvxzzjbdb@|+>Rt|b0w=zm8I6EaPv58=aYaYaSa<7kbKtFaFaDaK7M*0b29vwcbW+Ihu9IhdbBwtb0\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"{XaJvQaYa.bxwSa@u*bXaDqDa=qUm\\\"\\\",2):f(\\\"\\\"}qc.jb9bdbVaxb\\\"\\\",2):f(\\\"\\\"{*\\\"\\\",2):f(\\\"\\\"}bJdDqAas2ubTtRtOahbab<0Aawbiz6bcz+ex:wxkq*biim6\\\"\\\",2):f(\\\"\\\"{.jvYp?|C0>;cb6bZagbg,d+usss0w0:\\\"\\\",2):f(\\\"\\\"{=rpn,wp1=mz\\\"\\\",2):f(\\\"\\\"{bVa9bDa\\\"\\\",2):f(\\\"\\\"{bi/7bX2Ta7blw7wgbn,ef@|grvb6bDaFjSaPa0kjb=a2p2bix\\\"\\\",2):f(\\\"\\\"{8p*tx0,+hk;EaR-lbQaP<@qmb.bVa2<b.K5a-M8;6fkR1S1T:YaErWaAaP-+:H|o2X24bjb6bH5Zajbeb4bq.Ea/b?7x/l|QaEaj/:\\\"\\\",2):f(\\\"\\\"}vbDqPa6<o,z9Sav/M,djO4X-EaabdjX5Q-@ambnt.-0b?\\\"\\\",2):f(\\\"\\\"}lbubfbPakbUqcbAa:u-bTwr2xby,0babHyf99+mbdb*|w*u*UkBrhbBa-q/besCwf;zbcbcbgbSvCaubH5xvmb|;iq=xm\\\"\\\",2):f(\\\"\\\"}A5wbTrxxQa@a|4Tu@,kb0bSvUaM,lbXa3t+c>aBxcbabW+BaamOaM:\\\"\\\",2):f(\\\"\\\"}qes/z0sJ-Kp?a;ufbp:tbVaH5Xa-z68|b0p5bfbLuVak*i*<7@a\\\"\\\",2):f(\\\"\\\"}bIwF6ubj*0,ab6bXon|Z9a-R:Q"));
$write("%s",("1I8-b?aCt>jub4.2b-+wbGpes<\\\"\\\",2):f(\\\"\\\"}7bYai\\\"\\\",2):f(\\\"\\\"{kvI03j4bfpkwfsft-+s6\\\"\\\",2):f(\\\"\\\"{qd5*b4b*2wu*b3bkbzbvbTaOa.bEo<aG8guX--bFa0b,3+\\\"\\\",2):f(\\\"\\\"}hb-bJ,PaYaRud50*.*;j0s/\\\"\\\",2):f(\\\"\\\"}4yjbpq9pXafsD5vb>aybv3|/Va43Wa|.Qau|s|/bUalxw7A\\\"\\\",2):f(\\\"\\\"}Qa293vDqQ7mb3zUa-bB0x,B0L\\\"\\\",2):f(\\\"\\\"}@a9bAs,dS*5b>aar>apuL*0bQ.Ua6b|bub/v?o-bkbDwU\\\"\\\",2):f(\\\"\\\"}wsyb4b2h|bRa,b>aA/y+vyc8d9NaPa=v6jlwX0?11bFa4izbYxI*IpC\\\"\\\",2):f(\\\"\\\"{f+@akbL1I74-V|5s@au\\\"\\\",2):f(\\\"\\\"}-yd|8/:6v486ybZau\\\"\\\",2):f(\\\"\\\"{,b2bo|dbxb,+Ca3bdjTaSa/bT6ebAambcbhbd1tbWabvnxmb57c727yb*bDakbjy9be82+-b9bybC6,b.bq7hbq.5b=5Na+bJn:,6b\\\"\\\",2):f(\\\"\\\"}b,d5b1bOa=ti\\\"\\\",2):f(\\\"\\\"{wbNa>7R+>a?mEaqw\\\"\\\",2):f(\\\"\\\"{bHrs+UovbSvYajyubb4ms=x0bJnFapp@+|pUa1b8b+b.4N+xb/0Ra2s361640ub-,7bF\\\"\\\",2):f(\\\"\\\"{y,2z=a9bXacb>h"));
$write("%s",("6q9sC6h1Uaib+bCrf+fg.32bEag3hbI6ydK6Q.Sz=axbDc26RiPwub2g1-1beclxVacbfb>at0fsAaE\\\"\\\",2):f(\\\"\\\"{>a8s3j=qUa.uBa6b.bC-FaZa/uubtbe\\\"\\\",2):f(\\\"\\\"{|mS18*-y6*O1Ravb@pDc=aQaebxxPzWaxbcby,j,cb7o>-?aRambDqN|Xaf/,babKy:|dbDqYa9xibbbOoKtdrEaCawt6bXaL-h1Va3bTaZalbu*jymb8bebv|4bRt@a3blb8bWaVaGaK|R\\\"\\\",2):f(\\\"\\\"}QqO*gb44etIwYaDq5biblbo|\\\"\\\",2):f(\\\"\\\"{xFutbYambzbTaa\\\"\\\",2):f(\\\"\\\"}P0lqGpeyXa7bOavbtpn5-bAaJq4bRah1|b\\\"\\\",2):f(\\\"\\\"{45b/syvebPtebzkyu4bdptbUabb\\\"\\\",2):f(\\\"\\\"{bXawbUoDqCp3bn\\\"\\\",2):f(\\\"\\\"{4bP|I+1b?+xs//Aa@aT-\\\"\\\",2):f(\\\"\\\"{bAa2bk2v,qsjy.bkz@37b?\\\"\\\",2):f(\\\"\\\"}cyYa01xbz4nuWaws:\\\"\\\",2):f(\\\"\\\"}<tlb.bibYa\\\"\\\",2):f(\\\"\\\"{bdbfbCtvbM|=ayyz,\\\"\\\",2):f(\\\"\\\"}bwb?aH3-yOss4e|d-U17/N1:\\\"\\\",2):f(\\\"\\\"}@aab=rVxtuUa/bDqNaOaAaPabyTaPamvuyubmb/ktydbss1bit=-6bo1FretvbebQacb238zBxBacb>"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}ubgb7bswFae3wbPazb|36bbcQaErCaFgibL|Cqgb\\\"\\\",2):f(\\\"\\\"}b9ujbXaNoOax3\\\"\\\",2):f(\\\"\\\"}bRaCafb/bfbgs*bmbetR+Sr.bWa0s.0E+3b\\\"\\\",2):f(\\\"\\\"{bFaybEaWaabDqzbH2F2t-Qa9b>0B,2bTa709bbbp\\\"\\\",2):f(\\\"\\\"}cb6u6oVambdvBafb9b*b?aCxWazt2zYa-rwh*b\\\"\\\",2):f(\\\"\\\"}b/bv/kb=abbTaYoAa\\\"\\\",2):f(\\\"\\\"}bW\\\"\\\",2):f(\\\"\\\"}N\\\"\\\",2):f(\\\"\\\"{ybUaAaNa6stbgsO,.wwhf\\\"\\\",2):f(\\\"\\\"}7bgbTa4bCrabnx0b3\\\"\\\",2):f(\\\"\\\"}/buw4b6b2b>oj*dbdxb2JdSrQ.E1C1|bA1Fz|m-yUpb-;/Z,-yWp=/Cau\\\"\\\",2):f(\\\"\\\"}yb0bhbDqDqg+Na8b\\\"\\\",2):f(\\\"\\\"{bX.cmNaWr2b9g>,Mq.so1@\\\"\\\",2):f(\\\"\\\"{6bxbgbYhj1h1nxGx/bab6qgb|flb<aez<afb=a>uF*kbYa>hYaRoAaoxp\\\"\\\",2):f(\\\"\\\"{Paj.h.L\\\"\\\",2):f(\\\"\\\"{zbw01b<aQ0Yaewab<aFawb6bj,wbOaDqcbI+A-vblb,bUqXx4x7-UqtvZaVvCa2p3bW\\\"\\\",2):f(\\\"\\\"{ibjbgbXz.bYalbabE\\\"\\\",2):f(\\\"\\\"{8bwbN\\\"\\\",2):f(\\\"\\\"{1bWa+p0b"));
$write("%s",("ibqw:oDuvbOaixhz0b?tWafbZa1bYh<s>aX+ib>aD+.++dj0Fa2bZrfbIpDqfbvb+bPabbhuBaJoazbbRalbBaVmp/CojbBa?aW+d/FaYa3jt+OaWa4zOa4z|.x/X-7b/bi/VpGvV,Y,9/W,h|c-7*FccbVal/q/EtRaVabjEa6r9b0b.r4bvb0b-.Ealbgb+bDqF.mb=aSaH\\\"\\\",2):f(\\\"\\\"{VaBa@aAaVaUai-X-yygbdb?au*ebn-s|?ayz\\\"\\\",2):f(\\\"\\\"{.,-Dq>a3bCaRaAaOa@a2bibH-i.DaVaCkHy-.=aVar.=aPaSa8blbSaSa=a+b?aT-mbXaUa+qp-.b@aX-=aItOaXa?vRa8b0hRa>aEaAa5t+bU->aSa2\\\"\\\",2):f(\\\"\\\"{ybyyCz?m3qmbab/uhb\\\"\\\",2):f(\\\"\\\"}q@aWaWaTa<aEa.bRa>-@aSa?aSaVaSaAa7bDqTa:otbabN|kbmb+b6z/sabCaxbBoAaeb\\\"\\\",2):f(\\\"\\\"}bib0bhxdzFg7bWa3bibebCaPa@oTz@a7bcbyb>a+bcu\\\"\\\",2):f(\\\"\\\"{b,b5|0p@o6b*bkbSa\\\"\\\",2):f(\\\"\\\"{bU\\\"\\\",2):f(\\\"\\\"}Va?awb/++u6p>a7bB\\\"\\\",2):f(\\\"\\\"}=avu|ma-TsjkX,Qswi9*:*4*vbibWalbgsbblbPa7b=aCpzbhbUaOa+b<,4b+b*bU|htC*2b*b>aOa-bm+,bzbo|.bKybbUaa,Ra;pZr8bQ"));
$write("%s",("+O+UaFaarebwbRaNakwlbmbNaabaq0|UambOadbQa3b,bX|dvRaKt?azv>j4\\\"\\\",2):f(\\\"\\\"{dbHrvufpSalbbqV|9+/b+p@awbEaXaOa9zLuOamb9f2+zb0+bukbmzvbWa4b\\\"\\\",2):f(\\\"\\\"}*ubWa>j8b3bRiwba\\\"\\\",2):f(\\\"\\\"}PawuCadv+bRacbkbfbWtq+x+Bqu\\\"\\\",2):f(\\\"\\\"{SoUaPaHsN\\\"\\\",2):f(\\\"\\\"{k+?a4bzb@a?aNx*bC*zb<aUvTz-bOa0b,lii?*lb-bku@a-bfbn*/wibAaiiQlkzYa9bn\\\"\\\",2):f(\\\"\\\"}Kpm|Catb0b2b<aLpC\\\"\\\",2):f(\\\"\\\"{OaXy*bDq0b/\\\"\\\",2):f(\\\"\\\"{OiPa-yVs2yPnVpDvyif|vqQa*\\\"\\\",2):f(\\\"\\\"{|bVaGgesbb2p;uDa8babYa7barxbAalbFas\\\"\\\",2):f(\\\"\\\"{+bTaYaZo<aYa*b7stbebgu6bPc>a5bkbFgEtOuwb2i@aXalbyb\\\"\\\",2):f(\\\"\\\"}b9bO\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}b=|lyJohbXacxibZaNa2tbz-pPvDaDag\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bibYzfbQa8bZ\\\"\\\",2):f(\\\"\\\"{iq+pzb=aix=a7bDazvtbdrOaFa3bAq|bsuPatbzb8b=akbgbuf,bv|hzZa=aub3bFa-bhb>a>\\\"\\\",2):f(\\\"\\\"{@qkb/b\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{b9uEo,bcmfw*b+b,bOaVi\\\"\\\",2):f(\\\"\\\"{pPax|ZaibSaubii.tpzUaTaAiUtB|gbgv\\\"\\\",2):f(\\\"\\\"{bUtibiv7b1beby\\\"\\\",2):f(\\\"\\\"{+bijmbWa?aub\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{=xDq/veb|b2bcbTavbvb<o2gixebYaubSxbbbb-bbb5v*bnvQa0b/bSambbbyi0y1yc|Psgk/y8bbb8bkbcxy\\\"\\\",2):f(\\\"\\\"{Ea+b>s*b,byjvbUaN~2aeg-b?p9babNa-ttbPaKjjb/b.bmbsx+d4\\\"\\\",2):f(\\\"\\\"{Lo<abbarjbZa,b|rab7p,b*b/b5bvySawb|xzx4b@z6xebtbtuxbkbNa4bZaQaHsjb=zhb0bUazb\\\"\\\",2):f(\\\"\\\"}btb9bZaxsubabzbQajb\\\"\\\",2):f(\\\"\\\"{b4bhb6pxbyzDa0b0bAaababLi*b|bxy2bdzbz9zdb/b4bXaSacbOamz2qdbabTa3bubPadbYaXa0bkbOa/bnpVaxv/bAaVt4blb0bTuAa.bnpUo,b8bxyzb*xtbBaOajb>awxzbgbib3btt2bAatbbb=aOagpdb4bmbii<vAaTaFi7b9bcb8b-sqxEaVtmbibBaWakbZa5babgwPa@u.b=xgtDu3bXkbbXa<a1bVayi+y,ywi*yIbFvRnbkEvhb9b4b9xAa=xXx-bDq-bvwabXx6pou>jBaCa=xvbBa=x/b7bXaPa?"));
$write("%s",("a9bjbNa\\\"\\\",2):f(\\\"\\\"}bNa/wub7b;tkbLpeb5xGaJx1xJqiifrRatbcbibXkyb-b3b6p9b9btbgbLt1bdb8b7qbb.bXkDq+b6b,x-xDqiu,bwtRaXaNa?qxbXakb|bibgb2qNadb-bmbBa9uNaFavb8tCadb*bAa2slb3bXa\\\"\\\",2):f(\\\"\\\"{b?aJn6b\\\"\\\",2):f(\\\"\\\"{f\\\"\\\",2):f(\\\"\\\"}bow7bBa9b7b0b1bfb4b>a|bXa5b/bgb1btbOa4bPacb*pBsmbjbPqfbhbOaPaRawbbbvb*bgpCaQa1bPa0b\\\"\\\",2):f(\\\"\\\"{bgpPvCa*bwbZaXaQa|b\\\"\\\",2):f(\\\"\\\"{b-bZa7b.b6qdbbbjbEakb+bUacb5bdr<atb\\\"\\\",2):f(\\\"\\\"{b/bcb6smrIr7uebEa?aDqwb\\\"\\\",2):f(\\\"\\\"{b@t7bZa0bXa\\\"\\\",2):f(\\\"\\\"}b+b=u6bTr|mwiUsBvQpVpNsdbBalb\\\"\\\",2):f(\\\"\\\"}bDqmbwbYa3bXuublrls8r=a6bfb6oBagbxbKugbjbbbOaeb.iXaDa|bDa1bXa,bxjeb5bEaYaCa8b.bTaQa*bEaubzb/bhhRa/bkp8tNanu1hGukbVtZaybecZaKj>j/b=anuNayuzbzbitcbjbXkabibhbYabb.jYaabvbSaYaxb7bRolbOacbKpBa5bcb\\\"\\\",2):f(\\\"\\\"{bOalbbbQaCaOawbMo5bYacb*bgbKp,b=aCayb@aOa3bbq"));
$write("%s",("6bkbFa?a/b-bRaUajbab\\\"\\\",2):f(\\\"\\\"{bypmbgb*b8b0bdb\\\"\\\",2):f(\\\"\\\"}bPalbDq\\\"\\\",2):f(\\\"\\\"{bWa0bMhOaZp1bSaabQa?aZs4idbgb,b6bTaab4bWa|bDqSa6b7bFaibEa4bDqyblbTagbZb.rWa8oFaqsos5bwbCaDqib/bibQa7rkbWa,bFaeb1b,bWaCaeb3j?ayb\\\"\\\",2):f(\\\"\\\"{pcsSazbVpYnRsWnjmQnRpVpPpNp.rjbXrVrTrlb9bPrNrLrGaJr@a/bPaTazbab@a9rwbwb7bNa/blblb+bXaabwbmbubvb\\\"\\\",2):f(\\\"\\\"{b7bjbybjdhbYpWaEaDqfhubDq\\\"\\\",2):f(\\\"\\\"}bdb6bdbwb2bXaCahb8bgbablb\\\"\\\",2):f(\\\"\\\"{bkbybfg>aeb|p1b+b-b\\\"\\\",2):f(\\\"\\\"{b1bkb9b.b?aebeb2bUaiiprRaBa*bSaTa=r>aNaic=avbcblb5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaSa<aubgp9bzbjbRazb2bScebkrQaWaDqVaCacb\\\"\\\",2):f(\\\"\\\"}b7bfb-b1qDq7bVatb.b7b2b0bHqFqDq*bZa\\\"\\\",2):f(\\\"\\\"}bUavb@aoq+d\\\"\\\",2):f(\\\"\\\"{b-q=qdbSa\\\"\\\",2):f(\\\"\\\"}bkbdbib4b,b,b7bdb0bPa,bAaxbGavp,blbUaQa>aib,bebVahp\\\"\\\",2):f(\\\"\\\"{kWaBaFa+bSa3b3bU"));
$write("%s",("a4b\\\"\\\",2):f(\\\"\\\"{bebmb3bDaYpmbApzb?e;p*bBambPa8ojbFaPaCambFa>aTafbibOa\\\"\\\",2):f(\\\"\\\"}phb6b0b8bPa|bAaFa|bVp\\\"\\\",2):f(\\\"\\\"}mSpOpzmXnUn|m|m3aVnmb0bcbMhjbkbPa4b+phbNaBaDalb4bBaibwbhbvbkbvb2hZakbibnpkb?a+bfbwb5bXabbCajbTa\\\"\\\",2):f(\\\"\\\"{b2bfbYaiiqb4bDaYadbvbzbDaFa/bjb5bebhpjbcbwb,hDaBftbDavbdbPaEa+dBazbZa.b-beblbzb,bNa7bvbCaEahb<aCabb*b7b?aQaub*bWaQagbSa,bEa7b6bAaEaBm\\\"\\\",2):f(\\\"\\\"{oMmloeocoXftnzovo;alolnjncoko3mpo-blosnCa2mCnwbic8aGn=n>mfoEa2n\\\"\\\",2):f(\\\"\\\"}nan-aznWmUm|mbkSn\\\"\\\",2):f(\\\"\\\"{mOn9ayilmmmyikm|m/b\\\"\\\",2):f(\\\"\\\"{f-a9hub>h|e4n7nAaqn;n1m9aEaOatnCaMm0n6k:a,n=aEmYmcn4mqnCmgnhl<a-btnxnDmtnFm2mpnsnAa:aCa8amn>aEm=mLmGm8mOmAa?a>aDm|eXmzb5mIm6m@mBa2m<m:m*bvbtb/b-aJdHd+mHm?mDmBmSe|e;mAm?aAa-a1m8a7m5mFa@a2m\\\"\\\",2):f(\\\"\\\"{b0mHa.m9a|e/mxb8a+e-a1beg+mYl8arb8aXf|m"));
$write("%s",("4aymnjdknm?a5hPkPjkk7ejjhjUjbkimikikekyihkRlhj6b-a+czbxbubHaqb6aqb2i3i1i5aqbebCi,bAfzb.bKfnb|fldiiZgXg\\\"\\\",2):f(\\\"\\\"{gag|hSjwlthultcBaljzlHk.lDkBawkNhIg1iwbPfnkOk9k?aBk6e9hrb3b?k?a<i<kuhEk@aCalj2b3b4iUf?j8f6k-bxk@a3aKa\\\"\\\",2):f(\\\"\\\"{b;a3gwbccIa3b1bGj,b|b0auhmhuhRjlknj@alj.bri?a=kmk9i:kBa>aljybPc5kmhBhqj4hOjDa3a;d+cKf\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{gsbubwbii-aykwk:a;btk1b0b-b3a?a3a7b-aii.a:b:b,b?arjQjpjNj4avifkfkckNjwiak-fxikj5eijmdViRfmh\\\"\\\",2):f(\\\"\\\"}h;iPakiojmj9hwb+b-aPc;j/b8b1bPcxb;aUf-b:fZapg|b.b5b-a3j+i3bWfvb|bIg4ipgfg3bgf;a<b:b3b-a8bIg,bxb2b2btb;amhUh:iUh3a>a3a5aGhYixbWiUiabVaTaRaOaHa6eEfMhFfjb-agbebbbcbZaVa-abbVaEf-aZabbebSaHa@g-a2hhbQabbZamh4hjiWh\\\"\\\",2):f(\\\"\\\"}hQgnb-a2i/b3b4b.bHa8byb2b2gtbWfxb5bufid.gui/ath4a-afgdgMaFa=aUh-bWhBhAhGa+bJdPh9a/b5a|fC"));
$write("%s",("c8g-bPaBaobBhHfMa9aMaIa5axb3b.b4b0bxbzb-btbegmhkg4hGaMbHg2bzb;azbLfccJa7bmhth\\\"\\\",2):f(\\\"\\\"}hCdYaOaVafbVaibNa=auhuh?a;aSgVaNaUa.gthkgvbpbEa*c7bcd?aDa>anbJdubSczbPfIcQgyfwfuf2bsfNd3bHa?e-a-fZf:aIa+c9f:avbldub4bcb-b3ggc0gHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bdgfb/akgzgtbxcRf?a1akg-a6a5bhg>azd:a,cNahgwb.b;b>aagob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a,fPcFf/b:b6aKa6e1b4eIa8btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8a\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"LdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bld"));
$write("%s",("jd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})821(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,23^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Z3(yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalc\\\"\\\",2):f(\\\"\\\"{4sfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajn4bdateg@"));
$write("%s",("3doa2 kcats timil.v3dga]; V);R4aC3ecaL[c5aY4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.=5koa(=:s;0=:c=:i;)\\\"\\\",2):f(\\\"\\\"}4ajaerudecorp03gqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{/3bianoitcnufU6|sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fla\\\"\\\",2):f(\\\"\\\"})36(f\\\"\\\",2):f(\\\"\\\"{#,43z3mba7D3a835oa(etirw.z;)tuo.N7aba(66b~auptuOPIZG.piz.litu.avaj wen=zv4,ka93623(f\\\"\\\",2):f(\\\"\\\"{#t:355aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/n45da*6 L46ea1312~47\\\"\\\",2):f(\\\"\\\"{47fa41310?35Y9[83;M4dma"));
$write("%s",("(amirpmi oic$4[83jma++]371[]591[j55pani;RQ omtiroglaH35va;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})867z3a(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632|4,ea5526s@ajatnirP.tmfR@cfacnuf;P35datmf<36garopmi;PBagagakcapL3,ea3608#5dbapo5-?3cba-934jatnirp tesw:-ca69;;afantnirA5-ja9191(f\\\"\\\",2):f(\\\"\\\"{#f>31ca59$6awa,s(llAetirW;)(resUtxeT4Daca=:|5-ca38kAafanirp =33daS C;3-S=bca&(v43ba U4[U4qiaRQ margo#4/B3bjaS D : ; R*451B[83jL44qa. EPYT B C : ; A:5[83Cka)*,*(ETIRWD56haA B : ;A34ba [2c^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\","));
$write("%s",("9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'47ia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohce-A.ja(f\\\"\\\",2):f(\\\"\\\"{#(stupfEcdatniF3tca01z3sea%%%%:3[z3ipaparwyyon noitpoG3uw3Gca(n^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Csba1p@a\\\"\\\",2):f(\\\"\\\"}7qba5nIa\\\"\\\",2):f(\\\"\\\"{aetirwf:oin\\\"\\\",2):f(\\\"\\\"})8(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3c*8nka(f\\\"\\\",2):f(\\\"\\\"{# cnirpOAoc8dma.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\"));
$write("%s",("\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[06x#3cy4a\\\"\\\",2):f(\\\"\\\"}8cpadiov;oidts.dts vIaz5nV3d\\\"\\\",2):f(\\\"\\\"{3kkaenil-etirw64dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\"));
$write("%s",("\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^I<c/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qes"));
$write("%s",("od(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\"));
$write("%s",("\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\"));
$write("%s",("\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4)"));
$write("%s",(":f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.o"));
$write("%s",("ut.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\"));
$write("%s",("\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule