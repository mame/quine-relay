module QR;initial begin $write("%s",("let s=(\"Module QR\\n\")\nput=s\nprint\nlet s=(\"Sub Main()\\n\")\nput=s\nprint\nlet s=(\"Dim c,n:Dim s As Object=System.Console.OpenStandardOutput():Dim t()As Short={26,34,86,127,148,158,200}:For Each d in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import :wasi_snapshot_preview1: :fd_write: (func(param i32 i32 i32 i32)(result i32)))(memory(export :memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export :_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(d):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(6"));
$write("%s",("35555.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n=(c>124)*(8*c-41016):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^"));
$write("%s",("nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^6"));
$write("%s",("3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3dba;+3nna3(f\\\"\\\",2):f(\\\"\\\"{#qp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]#3sv3r23)ga7(f\\\"\\\",2):f(\\\"\\\"{#.33)ca51h4-ba1S4w23F?7d33&r7u53sda,4353.ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCL4/v4+ja36(f\\\"\\\",2):f(\\\"\\\"{#DNEm4[m4ada. A~5[p4deaPOTSn4[#5e~5[o4boaRQ margorp dnex4[x4abaS*5[m4c2<[ca91j4[j4eba&%6[l4bgaS POOL)<[:7dba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'j4[j4[j4gda&,)(6[?>cga. TNUO<7[s4bfa(rahcg:[(5dgaB OD 0B>[t4cca&,,<[,<aca)A36[;=e6=[.6cqaEUNITNOC      01z4[c9c,5[W8dK7[aGeeaRC .p4[p4aka,1=I 01 ODt4[TKecaPUq4[/I[6<hva;TIUQ;)s(maertSesolC;^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Ye%4Rra744(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})215>5[qa^32^\\\"\\\",2):f(\\\"\\\"})959(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})420pY4d8,ba8AAbg8[da304zY[O7bda218lK[wL[j4ldamif+6[ga)91361\\\"\\\",2):f(\\\"\\\"}5[,6[j4lbat(6[(6c%a315133A71/129@31916G21661421553/04[04cva%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})48\\\"\\\",2):f(\\\"\\\"{3bhaj:+1 j@34[34cbawm4[m4cl4[l4cbaWm4[m4cba\\\"\\\",2):f(\\\"\\\"{m4[m4cva)(esolc.z;)][etyb sa)t=[#>[j4[<6hea3289m4[x5[j4lba,l4[w5[j4hla!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~~v4[%5[j4hea(rt.o4[z5[j4hba)A7dda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};l3efa~~dneo3hra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a63j$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||13jda#-<q3jda||i)3mhaBUS1,ODs4qka)3/4%%%%i(N4cx5kU4xPa2=:/t"));
$write("%s",(";2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*45oi5vv3jd7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/rZa|atnirP/oi/avaj lautrivekovniJ3d.4j[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);24122<i;(rof;n)rahc(+K4r[2k*3&oa=]n[c);621<n++r4aqa0=q,0=n,0=i tni;N3&kc1m4asdRbQehmxfvfamRf<bedPdck\\\"\\\",2):f(\\\"\\\"}b;agb-a|dzdxdRfGb8aqeRdYd5a\\\"\\\",2):f(\\\"\\\"{b2bGi;agb-epb>a8adewj>aJaRaAdteFbaeIfOa5aacDg-b6f9apH4aLa7a;a4a<aPhnnkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9apH5d6cRbC3gUc-f/aof0fRfCa>a5a4m.b2e6aRa;dNaxbog*+Gh;aTapc4aLcEeyiof6amc<byg-fFmsbv"));
$write("%s",("h@CWfybxcxc>aGaUeAa2a6a\\\"\\\",2):f(\\\"\\\"}g7a6a@a\\\"\\\",2):f(\\\"\\\"{g:a?aMbKaKa6a?e:a0A2a|gZfMbbgli>a:b1a-glnUf\\\"\\\",2):f(\\\"\\\"{bHaucMzS\\\"\\\",2):f(\\\"\\\"{pzX5pzEc7>JaMa\\\"\\\",2):f(\\\"\\\"}bJae1Ec-bJaJaP\\\"\\\",2):f(\\\"\\\"}JaMdJa8bO=;a8basKa8bas+4fkj9Oac=TG9bKa8bSaA,Ta8bC.as8bTGJ=JaLaJa8bC.Nah4c\\\"\\\",2):f(\\\"\\\"}a8bNa-9TG:b+bLzfkLzfk\\\"\\\",2):f(\\\"\\\"}bJaHaJa93c/aHaJaFdmC;a8bSaUa:aUa:aO=viSfQfNm4a81sbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'maviDa-a|bv+-a<6asal+Ue>a/j\\\"\\\",2):f(\\\"\\\"{gKaKa|gZfz6cgaagHkkg~6esasbvh*b-a/bxcHa|fDle3c0c\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{gph\\\"\\\",2):f(\\\"\\\"{gvg1a-g\\\"\\\",2):f(\\\"\\\"{b"));
$write("%s",("HaDlRf-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?a\\\"\\\",2):f(\\\"\\\"{gJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1a-g0iDlxcpb7anb2b:b\\\"\\\",2):f(\\\"\\\"{g2f7k@d-aIfVkxcHalgjghgal-aUf0ixiRf-f-gSf|fDlzeSgxiHaTk;a/aDh<b+hWh<apb/aDhWhnb<a,H:b\\\"\\\",2):f(\\\"\\\"{g/aDh-f-g+gFa,i|b1ali3b:b\\\"\\\",2):f(\\\"\\\"{g9hHaDlHaUe-iCe|bxc3b0a:b\\\"\\\",2):f(\\\"\\\"{gIa|bzeJa|c5buaQbxi<b=a-aAn*c3bxdUem3aea|b9ai3efb2bMa7arh|bphnhlhjh9apbqhohmhkhKcdc/bPcgfvfOhJh7aEa|b.l,lMaAn*cEc,dJa>a2aIfUjMgMaAn|b<i+cbi6a13kWaxd\\\"\\\",2):f(\\\"\\\"{,vb8g/aDh=apiJ7-cJ7OakbA5=xpi0k6a7b5aTkRfwbXjUe2b5a9g:jmPhcloOiOinq0c/bxd;a<hJj^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'?aea6a2bL>"));
$write("%s",("e\\\"\\\",2):f(\\\"\\\"}czC5M6a-o2a5axk2I\\\"\\\",2):f(\\\"\\\"}gEhgl\\\"\\\",2):f(\\\"\\\"}uOi6aUh9mHa1dmdLhRfNl7mHa:eNl7myk;almQaabRaRf\\\"\\\",2):f(\\\"\\\"}G<b3bxd6aIh:l5a*j7vkixb9iacPa;a9jccI?pbubld1bZb\\\"\\\",2):f(\\\"\\\"{VnbpgPjNjEc,d0kfl6m<b<b<b=k:b3k<b<b,cBk?k7b-bBkEa<o3bDdzlMi9a7b6g-a5b7|,cBk=a9a7bubxbs3e33eca:k33eea.b8fE3c33ifaJb7bd^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3fna2lQHBa>a9a7bw-3dmakiolKj9l,cBki3a?akn8|fh,cBksbHa\\\"\\\",2):f(\\\"\\\"}gmkMlkgKlMk;kCaLi6a0kflXkik6a6lWlPkUlxl<bzeWCc93gea1lLi+3edbm4A8tW0c4mqk2m0kfl?l=l3a6a<bki>jD*\\\"\\\",2):f(\\\"\\\"{S5MyS3M2a2a\\\"\\\",2):f(\\\"\\\"}GVkPl0iwbXjRf@a>anc:e7b5aWf=aKc"));
$write("%s",("Cusl5a,bJa6a/Aa%aub9h5aUgwbXjHa:e-b9a9b9adlVkyg>am3ayaXJVkyg@a>a:a|b9a0b9a@a>asCa?a>e|bPg9bJa0bVkyg-b9adl9aL4Ja9bVknbJa6a|b5a,bRf:e-b5acotb-a,<a&acwA8tWvi\\\"\\\",2):f(\\\"\\\"}Gyg8bAdGh-a\\\"\\\",2):f(\\\"\\\"}G?Cbb-a\\\"\\\",2):f(\\\"\\\"}Gyg7s3hea\\\"\\\",2):f(\\\"\\\"}G?a*6cca.jr6a5a\\\"\\\",2):f(\\\"\\\"}GKcjE/bxd6a-b9a8b9a7bJcJayb>aTuki>aJa*c@dxc?b57o3a1a-bEmteUe@a>a<a2b5aDcw3:atcJaub5aEcxb@:,bmPVgC;aeaJlHlQ;aP:aka\\\"\\\",2):f(\\\"\\\"}G7esktjpkn8gyaTlRlpb;awbXjsm*k\\\"\\\",2):f(\\\"\\\"{UnYyUoYQ7a+avWA8tWFcjnumPnuo@m2n0o\\\"\\\",2):f(\\\"\\\"{o72uoSmqp6,Ra5693a8duAlYwbc2<tdbXaCz\\\"\\\",2):f(\\\"\\\"{beywE1@2CBaxXmQhxEt0|Daww|basGauSH@0pa*oGLoo\\\"\\\",2):f(\\\"\\\"}RaTa96Lo=,3b7vKUVxMsZo5bpuL?Sr\\\"\\\",2):f(\\\"\\\"{QBa\\\"\\\",2):f(\\\"\\\"{zhbrpGLPaDaib@afb>a1pkd4wXac?jbvbvp=aqpryHp@a\\\"\\\",2):f(\\\"\\\"}/g-,d3qerDa2sYaEa3+rC2b=atbEtzrOwzwojEE"));
$write("%s",("Zam\\\"\\\",2):f(\\\"\\\"}Dalb;FN|2Y6,tb4w177,bb/So\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}zY0Aa7b:5mbEaVx.bebm./1VK1\\\"\\\",2):f(\\\"\\\"}KIsMYaj3zsL-+buxSI/bRGx9eb-bmbtb>3m.NamCkbfF|;ki4;-qaPIN/+Ra56*?c:yT.qf-<6e&dy-Y,5u@;Y<olZ>db7-Et-xgEvM0\\\"\\\",2):f(\\\"\\\"{RL>a7\\\"\\\",2):f(\\\"\\\"{hB/45b<an,s<Qu-b+|3H\\\"\\\",2):f(\\\"\\\"{b57V21b*<7bc90VXa4*y0bpq+X*J/bb@<db,GxbdIjbq=|bSz3YVvs\\\"\\\",2):f(\\\"\\\"{Sa/xSatsyb*bmbbbDaufq+Saf*TTf*Ra?ZWaVazuZF0ljbub5yBaNaj7buS+Ya1wh9z*>/kbi*.*2tQukw*4YLmbEa++|+t,Y0v,Cq\\\"\\\",2):f(\\\"\\\"{d>aJuW2Qr7bkzOypv2bWafrJI.+b1y-mpus+tz8kbT5y.Pwz5XaT5VzdbiOVa6bE@p15urr8|3\\\"\\\",2):f(\\\"\\\"{fp.+ac.6e)c:wfpNvMoZFe;FVY5AaYaj:LX1bK,Yaj:P3S\\\"\\\",2):f(\\\"\\\"{0y.0Q/6Za91w8H=Cw.r3bZA66,FTIADajbbC@aYq\\\"\\\",2):f(\\\"\\\"{q6|7W<0BvgbEpLoh-wJDa@4U-n@,b?+w.0\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}qs@*T|TzTkhF4V-eA<:tTq"));
$write("%s",("+qTCpoTgpu+yZOaYqop6,jWDDjbp@C9eAb1Ggj=y*w*UwZov<1@Ms1@wbkh<\\\"\\\",2):f(\\\"\\\"{Eau*jb?n?v6bCao3a7a@SX9y-nGlb2bssw8,bsFNa1@BaRaLU1S/S2s.,oTsFKRy-u*Zan6e@blbdp2y6ZU0@PUqjSw.EpBqQadug;y-6,s\\\"\\\",2):f(\\\"\\\"}Zo3s1@SjURSajbQaS+KNkbaskiI,w.jXbZkiV+asHR1@5bap7Khb91AR1@0FUau\\\"\\\",2):f(\\\"\\\"}<R\\\"\\\",2):f(\\\"\\\"}4i0iVO-2b7bCa<\\\"\\\",2):f(\\\"\\\"{=ae\\\"\\\",2):f(\\\"\\\"}2b7bubDadsZo5bDajbDa7b.b1@m3aObErAaXakC7bubErM/gb08Jw3bGLfb9bEa,bhw\\\"\\\",2):f(\\\"\\\"}brgxb6b+S7bSnDa|bEaKIq3Fab>tby|u/Mz/sTa,J0bUukbXrjb/sd6hbnhPrPpgbPaLq+AEambDaOy\\\"\\\",2):f(\\\"\\\"{j|pg4QqT*;wN.H+EirSFaerwbKpn2yIOa<<F=Zaz*DacQ9f1c.4f*.4ZaeX7b0bSYJ|7W=a,b8bI;/tn/QUvb?Im*|,0z=aStlTLHEzQH6.iB<aFW@n.+pF0wvb?I\\\"\\\",2):f(\\\"\\\"}t;|RZvySl\\\"\\\",2):f(\\\"\\\"}L\\\"\\\",2):f(\\\"\\\"}BTaczazhb/rzpRJt-<?0<>|0<eyVKEa+?WaO|dNq?iA0RH-F;B+O|gb,\\\"\\\",2):f(\\\"\\\""));
$write("%s",("}b5bbF;mb4x6jz8us9/DagbJU2bzHojXausD-.d/bxbL6WaE+jb46h:EaF;ZM/bjIib/xtb9/s3akar\\\"\\\",2):f(\\\"\\\"}YaybcWWa~4g/a4=s=M0gbnx|b0h?a1h+<n\\\"\\\",2):f(\\\"\\\"}Nar>.t=pr4P3JT|bd@4z(6evdFa4=U6+d=p7tWTVa1yabr4P3m\\\"\\\",2):f(\\\"\\\"}2Sr4Br@rr=2uq+|\\\"\\\",2):f(\\\"\\\"{jb6+Hq2SnvM8ypq\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{blb;EkSb76nhpb>y7O*@2PQjJJ0iR\\\"\\\",2):f(\\\"\\\"{AjbNS|2*bT0s=abFaozYa@-1bBMO>0RAajwVU,bH;.\\\"\\\",2):f(\\\"\\\"{YL1-mpQ;G:c+@a|bNaetPPb>*FsM<KkbE8q+gb*+\\\"\\\",2):f(\\\"\\\"{ln.3z9vh81lMLCrNaxbU8VQxbabu\\\"\\\",2):f(\\\"\\\"}2bLUW@ZEj6T*MC+bFabi,bpHn,Nqyd/ZUkmxgW5x-Bg9Ar?xGOtbWPh9Ez8H1xibQpvb:j/bwb\\\"\\\",2):f(\\\"\\\"{b++\\\"\\\",2):f(\\\"\\\"{V~6e+dAL0JALOa\\\"\\\",2):f(\\\"\\\"}bK\\\"\\\",2):f(\\\"\\\"{k@*,sx54k@5bgb,pzc8biRib|bHd0o6b<acQDtB,.+2+:=Tt,biA3bw3:uCrS1ZaLBAE<K*u<sCphI915b?agbu\\\"\\\",2):f(\\\"\\\"}2bCao8u9bbCwh8tI,da\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{91V6\\\"\\\",2):f(\\\"\\\"{yiv<qa?nLh:Dac:<:Nrzb?aib+bybZ\\\"\\\",2):f(\\\"\\\"{r\\\"\\\",2):f(\\\"\\\"{Ua=SUH*b4=bb+4=Wd\\\"\\\",2):f(\\\"\\\"{ZaEIY0uIOa\\\"\\\",2):f(\\\"\\\"{b:-|DjuML7b7bab1,UFHj;\\\"\\\",2):f(\\\"\\\"{,b5X3?;r3gQ/CahKBatxeKcK*bPa.bEau4wbjwdbYB>awb-lAav6M|mjWaebzbwb003>@4EZ70Gaw+0;S;Fa6tL6PeAf~d7hymt-eK4wdb+Px@zbx:Pa1xt+RavbjbfH<a@z09z\\\"\\\",2):f(\\\"\\\"{0b,zMVf+d+YaPCd/MLCrX.J2cr<aUa-IYhki7st+I=mRj7FVRO<.kb+bO=JVFVUU,b7bQ3CUVabU|:s+lbq+1VDvmL+*\\\"\\\",2):f(\\\"\\\"}*\\\"\\\",2):f(\\\"\\\"{*\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"y*w*1u7HM|aEq,1qVPUpUwTSBawJL6G:rg8/o\\\"\\\",2):f(\\\"\\\"{0hzXY7SMZaFVYa4vmb1\\\"\\\",2):f(\\\"\\\"}7qJT7qKv?aq:*Scr/rRD5brrhrVzHsu0g1ib|bz>5gybXrtbUaSv\\\"\\\",2):f(\\\"\\\"{lSar6DaOa*1u*+cebmvdb\\\"\\\",2):f(\\\"\\\"}bCa@Dxbc:59sl<3PaDv*6etdpr7gv\\\"\\\",2):f(\\\"\\\"{W\\\"\\\",2):f(\\\"\\\"{wbDTZM\\\"\\\",2):f(\\\"\\\"}qhxzxDcNaKxs>b>gb5\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}ebr3a\\\"\\\",2):f(\\\"\\\"{:sn2yhRS:sn2.bpz?aPaaiubGp0w82-2+2\\\"\\\",2):f(\\\"\\\"}2?w\\\"\\\",2):f(\\\"\\\"}YQap,<aNaWuWa970-@rlbi@KfdbG>?fh2a-Y,C.V,4bk5Paq1Jxxu0zaiubldT0*DfsV+qY07++6bh2Zzn/n+2be\\\"\\\",2):f(\\\"\\\"}vbvbjbn+zb0wvzfsI,2bLEuf0wi\\\"\\\",2):f(\\\"\\\"}bb2LVaBRUpvb,|,tiR+v\\\"\\\",2):f(\\\"\\\"}b7bI|rx91,rmb8uY\\\"\\\",2):f(\\\"\\\"{8u4b5z1bG,kWGLtQjI\\\"\\\",2):f(\\\"\\\"}bju918b||Jdf3Kx\\\"\\\",2):f(\\\"\\\"},j1Dt.bm:Ccs7aca,b(6ebbdbW20wCRT6XrAu4be\\\"\\\",2):f(\\\"\\\"}vb9V\\\"\\\",2):f(\\\"\\\"}/W7U\\\"\\\",2):f(\\\"\\\"}jstUn22|++Z\\\"\\\",2):f(\\\"\\\"{3bISEamRl<dr4xEa7-=l9\\\"\\\",2):f(\\\"\\\"{jb?afb>aYLzESa6=|bT,N=H8xbr4c^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\"));
$write("%s",("\"\\\",4):f(\\\"\\\"'c@-4bA5Eas6d@Oa45\\\"\\\",2):f(\\\"\\\"}bz-7rWagF\\\"\\\",2):f(\\\"\\\"}bz-c5O>K6o,,prX3z|fll\\\"\\\",2):f(\\\"\\\"}bYrLu1b9\\\"\\\",2):f(\\\"\\\"{8b4bkb-bSaH;5bLsHu\\\"\\\",2):f(\\\"\\\"}bmd\\\"\\\",2):f(\\\"\\\"{-Ua7PjS5G/Btb.Xgb8>/bmUkp/1rXNor3@ClbG:tUrrhu\\\"\\\",2):f(\\\"\\\"}A\\\"\\\",2):f(\\\"\\\"}b1bLEy\\\"\\\",2):f(\\\"\\\"{FJ7bt\\\"\\\",2):f(\\\"\\\"}y*XrTGa7Y0:0<aUWhbdbTNib+bvbOalbEaf+iLM/LEMz.54b6bwFogtb?r\\\"\\\",2):f(\\\"\\\"{b+,Ps\\\"\\\",2):f(\\\"\\\"{i$Vgbb<8;Lwt@p3bO-gD@Dx6\\\"\\\",2):f(\\\"\\\"{7H;\\\"\\\",2):f(\\\"\\\"}bebfbrTmbtb46@;kb6BeLjbfw8u<aub>3Ba,bKjRa:8Sa.+<azbabp;Nap1/bCQNaq3a\\\"\\\",2):f(\\\"\\\"}cFak054ib.b@DDle\\\"\\\",2):f(\\\"\\\"}vb.MtbQ/q\\\"\\\",2):f(\\\"\\\"}dgJ0vbUp,bslc5U6zN2Y+\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}2V3?|KG2LlGZucbTa;3TauRasbp/tTMwb0,q3P.\\\"\\\",2):f(\\\"\\\"}bk+lRGLW>Ks?D<a@zvb@uz*\\\"\\\",2):f(\\\"\\\"{bM02b.M@zt1RSwsLsH@JyA0lR4z1hLhb\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}t-g\\\"\\\",2):f(\\\"\\\"}D>f;tb=aX9+.fbETWa:FO+hbXsR+L*Wanv:5y<Y27bHu*bxbabW@l:e<bjbk*1VlAvbvbwvkvb>kuiuI/gb+y9z0zLqupXr=l5sk054|bi.9\\\"\\\",2):f(\\\"\\\"{mb=a0pnBw>f><a1VlA3qXqFt?=fhCY0zXaWqi*@au|y;=Arvz;lp|bh6Ps\\\"\\\",2):f(\\\"\\\"{bz\\\"\\\",2):f(\\\"\\\"{fk5rMN2*JxwQ<qLHtQL6R>2*7bA+D:a:b<aH/2*;9Ht@iGEEa9b>\\\"\\\",2):f(\\\"\\\"{7Gabdt6bebDv/Bb>9bTaeRPmUi,bdM-BkiIm\\\"\\\",2):f(\\\"\\\"{V52:0.>2b\\\"\\\",2):f(\\\"\\\"}Y/yeQCz/42y\\\"\\\",2):f(\\\"\\\"}Yt,jbMofboyu;GEab.y0?XarDxb<aMo?=J>O=K.j>F<5=6b<a,5@7QaCpR8P,(6e>bR8P,Qa6,INRaJD/2P,Io0w5bA,3;.r3<jS8wg2kb\\\"\\\",2):f(\\\"\\\"{bt+Ra6bs16b7wxwos@WQ\\\"\\\",2):f(\\\"\\\"}RaLHx<Ca/b..|bebq\\\"\\\",2):f(\\\"\\\"}Q\\\"\\\",2):f(\\\"\\\"{TQYCFqEE@W>ib3NaQ\\\"\\\",2):f(\\\"\\\"}Ra8,k*YaCah;ozovY0Oa/uoyRL4HGiTQS5.brTPrz:X+%3aeawFfbu3a,blb?xg1W3XtTpRo5bUab7Uauqiboy|mg9cW..b7@zzdO-E68P:/U2I8GsjdY7ld"));
$write("%s",("+.*b\\\"\\\",2):f(\\\"\\\"}4rT4Has6Ux2@;p,YaV29bvxGakBH@2bki|L\\\"\\\",2):f(\\\"\\\"},sw>Y,>o\\\"\\\",2):f(\\\"\\\"{-Hqsg-n2l<h2psZ@g;cO4-szbVHbU=2p\\\"\\\",2):f(\\\"\\\"}Q6,?5b9\\\"\\\",2):f(\\\"\\\"{8b\\\"\\\",2):f(\\\"\\\"}P\\\"\\\",2):f(\\\"\\\"}bP\\\"\\\",2):f(\\\"\\\"}ms<a.49S|w2yLqx-q+dbTaq+x@9TQ|Ow3t*B\\\"\\\",2):f(\\\"\\\"{bo\\\"\\\",2):f(\\\"\\\"{Ra*bUa9w.bfbnwq+Cpx@9T0HCsbb9>7F1MFaWauwybxBEaj:\\\"\\\",2):f(\\\"\\\"{bA1*bztuwCa+BjJZsuS+rOa=<FDW2?aJvWr\\\"\\\",2):f(\\\"\\\"{Dn,+bIvA9U0/bzLZsuSGRt*CrR\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}sz:7|/bp*>aPCAYh7>YOs/+qs2b:wB7er.br\\\"\\\",2):f(\\\"\\\"{P5Auvbjb33aka.bss+b0V0pE3c+aGWA9hbvTHqPap*3w5b.b6b,w+b\\\"\\\",2):f(\\\"\\\"{p<:ax<:3\\\"\\\",2):f(\\\"\\\"{Xs*6eTb+BJyzb57SIdbVHEaUa<a*UA9xY8ulh7b0bEabb-u=p/*ki4;sMNxzbOakzZM3BbbF@lRg1Wqh2=a8w3Qx9g2kj2rEqRJH,-brTg1y1-GOP\\\"\\\",2):f(\\\"\\\"{.UwTp7b>YGakB\\\"\\\",2):f(\\\"\\\"{bO=\\\"\\\",2):f(\\\"\\\"{"));
$write("%s",("DXq2bEaa5-l9+lGZuwbj;LrK,6sNqebpHn,jb7bV?i3a5a\\\"\\\",2):f(\\\"\\\"}-Na:|x@d/Pa\\\"\\\",2):f(\\\"\\\"}bR.Nxd/PaVav0HIz@tPc:+2Y6-+VL0O5<KEWEaGaiV7bVLtU;whvX+jXlbeY7lgM/zeYWLb+bbxbBaVQ4v|-rRWuRa.4ybz@R\\\"\\\",2):f(\\\"\\\"{h-54F8mj,6e|dVv7r.bg:ybf+lRjw0s8buxdGJK6beT5b0?>\\\"\\\",2):f(\\\"\\\"{c:b\\\"\\\",2):f(\\\"\\\"}/+kiRFPCzbJKvf0va\\\"\\\",2):f(\\\"\\\"}2S4P=a8wd52b=1-BNaZskBg46:pzbbdG*tDux3OVhBYabkJAhbTac54PW0vbz\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{b.sQa*b0<hw8HhxNrC6Ba\\\"\\\",2):f(\\\"\\\"}bR?EkvvZ/y\\\"\\\",2):f(\\\"\\\"{-bN=Da++Va36A0Crp7tGNabxQxbZnJMvPs;wyI>7Ua*bfbSNy\\\"\\\",2):f(\\\"\\\"{f;7b25j,WVCpw3jbT66bCxw3>ads:9bd3qmFb+bbtb?sz-RawpbzusQa9yDahbquS+QuUu6|g-??xy?>Q\\\"\\\",2):f(\\\"\\\"}+*EGi<b@**2dbv1BaVaRre;6B=piz/xRL6b-.>aWqZ+LuuvdKScRagbL-mShbI2xykzt;t>a*xbGz;w-bf;@PTw>ajbZ4lb0bibbrgb8bH;Mh;w0=ebyw\\\"\\\",2):f(\\\"\\\"}=1\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"}XwCz0<f6|TAKC7TaT5h<dbfc>avMKWa<bxbGaL7s\\\"\\\",2):f(\\\"\\\"}>iXjYajvg.dbTax<WyfuZEq\\\"\\\",2):f(\\\"\\\"}O\\\"\\\",2):f(\\\"\\\"}UvQag=-pJdWwTH3Qkr>Euu:/h.sJ0<tQebRV0@<?z;zb|b,BB\\\"\\\",2):f(\\\"\\\"}>7bbg6;r5\\\"\\\",2):f(\\\"\\\"{vbMq8sbZEp2bt,AQk@F<KfMr0R2b7bmL/=mbTa?vCa3D6bspLNghbeb:04Hzx/x48Gp5baRmbeV9b6beb\\\"\\\",2):f(\\\"\\\"}4f*dMU\\\"\\\",2):f(\\\"\\\"}tHI;uK8br\\\"\\\",2):f(\\\"\\\"{D-H;pHUaq/Cp5gM/\\\"\\\",2):f(\\\"\\\"}YQa,b>aOa|uVH>|Ua,b?wb+AabH.2@fIEc1aQaUH=C=aSJ;v6b7+5b5b8@?+p1Aah=>aSzt-nvl^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3mja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(|a3891(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})4201(f\\\"\\\",2):f(\\\"\\\"{#)~4[~4b|abQa*4tZ+bxbkiSKO+TaK@:/h.6/q3c%b*-FaSaiR>s,:uu*-xb0bbbYa+yW|xb=W3bd*7rWM"));
$write("%s",("Oy3@t2Ea5b-bbr8bbqZI3TOoGGR8p*g4p,/@g@5yY-V1p1*-nx5btvqiab>aC@eNTaGG>sayy</8Va3OFf9aJrayLjC1-+j@*-nx2+lbEa,:uu?abHVajT5sepTagxnvNaLL\\\"\\\",2):f(\\\"\\\"{D@a^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5e@cAtQHTy>@Y2;3?xf.hAVzwyq\\\"\\\",2):f(\\\"\\\"}WY*DQ;5\\\"\\\",2):f(\\\"\\\"}?aOph8TQ8XH;bbd\\\"\\\",2):f(\\\"\\\"{mb9bpw59QpN/>a0bZy4b*?;9BDbSebPCCwaEI,=ptbg-ufohevXa|+-bxhRa1b@aFVRauboM@alb|+qu@a,YAzTB1z0|NaFV1\\\"\\\",2):f(\\\"\\\"}L66b>awbFaZH<.2b@a|+PxjbYaxbaiKqco7W,rLvf*Oo:\\\"\\\",2):f(\\\"\\\"}JC?td<\\\"\\\",2):f(\\\"\\\"}TbqN8/3zb:fO|b?0b3JDairGzXaX,D\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}be06fecYaZTxbhIhc*4i|t51bfX?2,bjbKJ9b?aOwL|="));
$write("%s",("ryb5bS;FaWa<aQaVag./*Mv.G|N09uRWMV?cbNaJTg.\\\"\\\",2):f(\\\"\\\"},+.GoUMUan/SL8,*bDaeb6bO,pznsm\\\"\\\",2):f(\\\"\\\"{Fa=*=a,GVaeJ:Q,26b8=NNu9\\\"\\\",2):f(\\\"\\\"}Yd\\\"\\\",2):f(\\\"\\\"{:;BrUMf;tZq+\\\"\\\",2):f(\\\"\\\"},bvDamL3yx:,G+|Ya/sxrq\\\"\\\",2):f(\\\"\\\"}HBb4ipbzbIS9b>a3>1ln6F8NaxbVaub0v>anDTDg61b:5v4w\\\"\\\",2):f(\\\"\\\"}7P7IKMq>|L,dKfz@IS\\\"\\\",2):f(\\\"\\\"}bCYTDg6O\\\"\\\",2):f(\\\"\\\"{QFDz1bT24wO3I\\\"\\\",2):f(\\\"\\\"{8bd3SYeb?223P4Z?g4.6e,d-=g;+b|:Ua0ANaTaUwL\\\"\\\",2):f(\\\"\\\"{ybU0>a?aSj6nvb>symwb5u+t\\\"\\\",2):f(\\\"\\\"}tsls6AVTa7bOagFTGEa-pJdmUuF\\\"\\\",2):f(\\\"\\\"}b8bDqeb.bNyR\\\"\\\",2):f(\\\"\\\"}W2bbl*D+QxnnogPQksL60JUFZaNqdbcba*>\\\"\\\",2):f(\\\"\\\"}D>PjGgPj54-bmb*DZa>a?a9\\\"\\\",2):f(\\\"\\\"{f/g4NC+,c9c5b5cbnwfrLTzv4bswdbcbn+QaldUF3<Cs?C*,,b8S/bwbu\\\"\\\",2):f(\\\"\\\"{+px:PaVav73.lbCYK7yx3QbrWa\\\"\\\",2):f(\\\"\\\"}bP,UUeQXsubapbzRD5bMC04Ua+p.b"));
$write("%s",("6bvqwJg4H+gQ4?wb.tY0L-ou5;Kveb+HZ*dJ+b,z46e%dQo9VpHUaPs|*FZeuXajb7b<aPa|mjbdbN5\\\"\\\",2):f(\\\"\\\"}*Zawplbg=nGQa>fWQuS\\\"\\\",2):f(\\\"\\\"}beQcbIvnzy0fbtb1wkCRa:6+bWLdbcbmx?a71FV5vdVvbKHnzy0JF9tR3eGcmp9NrUkWuGakB6bdyastIHn<*vbdbdq3L<:0LZa?=,bR8fbAP?PVaWahI/bfI+PRJYatw?>lJqpquGz5sVamb1kfh-8EIeA4=z\\\"\\\",2):f(\\\"\\\"{Aa/b6b4\\\"\\\",2):f(\\\"\\\"{0b?a;2RmOwcL8D??eLoySap\\\"\\\",2):f(\\\"\\\"{-p@4GaL7c*UBw=i6oJ8,,b/byt++6b?IEtSni3;\\\"\\\",2):f(\\\"\\\"}Np3Jwb63=fsatEIwZ*hU4UWChB9-*bK3efdtQ7bxuJwe\\\"\\\",2):f(\\\"\\\"}kzlb@0QF1|iwhcGOWu-8JpuFNNRa3QbrON0-0HmHev848,Ta2b7bSzO@,b58.V;P\\\"\\\",2):f(\\\"\\\"{bqu<adb6bEcvb-bubc.Sz|\\\"\\\",2):f(\\\"\\\"{M0,A2b\\\"\\\",2):f(\\\"\\\"{s1lL\\\"\\\",2):f(\\\"\\\"}0<Ps<aUau\\\"\\\",2):f(\\\"\\\"}A,Pa1\\\"\\\",2):f(\\\"\\\"{pSqp6,Ua5g5G=Sh/>aVxjbH+bbBA7\\\"\\\",2):f(\\\"\\\"{ufn<gv5\\\"\\\",2):f(\\\"\\\"}Scg6zbgEf>7l|I7llbW-@Ny;|"));
$write("%s",("-0b?a2bZ\\\"\\\",2):f(\\\"\\\"}ywhroJ3beb+.|b,UR+gblbQa6B.bn.eb6JzbtE*.|sfvJdfbbQJ>z/-bSa6B0h7H0h=agNi(bFcg6TuwbbbIoXqkQM87qyxgv5\\\"\\\",2):f(\\\"\\\"}gvKu3<v@WayxurRPScg6gvRPIsUz7bzbXq3b72cb8BXauKJrnJ+bx;OVJ>1zF71zF7Can/5Y@Yqp8b:Ufbe1Eabbydps4bxbe3avaT1yd\\\"\\\",2):f(\\\"\\\"}29g\\\"\\\",2):f(\\\"\\\"}29gybMzqr,p7\\\"\\\",2):f(\\\"\\\"{3b4bSaecOaoB/xyb\\\"\\\",2):f(\\\"\\\"{bBaWowzW\\\"\\\",2):f(\\\"\\\"{6b7\\\"\\\",2):f(\\\"\\\"{=\\\"\\\",2):f(\\\"\\\"{,Af*.+u9Zq4bf+PSF:RabbxXHquuCQCsqpfrybGiJC3urI/rzb\\\"\\\",2):f(\\\"\\\"{sEH,bTa0ba@=Shs=SIKVKvbzsYrm\\\"\\\",2):f(\\\"\\\"{KEKRr=.+2OkbBY6b4\\\"\\\",2):f(\\\"\\\"{WK?v\\\"\\\",2):f(\\\"\\\"{bO5Y9ecc\\\"\\\",2):f(\\\"\\\"{sy*Jh/bdbEaFf|YvBfbxy.Yjb<KrIf++Arjh/pROy-i\\\"\\\",2):f(\\\"\\\"{xCpM>@;:F8sab=0p1?a,d0,2bH;Uwmbkiq,RONavuGE@S+yWqtbKxjwhbEaJ2rTos/1qPgb:-zb1k5gNS433>IROPO5-xt>Ra9fhb7Kd0Ft0buf-CY9,bUaY2\\\"\\\",2):f(\\\"\\\"{"));
$write("%s",("DBY6b:U?=[NctbF<Kfvp6bebFa@7p1PaR0w3Oy58P4bbpHp1Wx-s<awbss2bRa=r/b/xj6xB2bxj=,mb*<5+E33uLy+b|w-95|FkP,lGrrwtlbJ0-bOqkb7l*6ewaDa7b\\\"\\\",2):f(\\\"\\\"{=8>\\\"\\\",2):f(\\\"\\\"{J>1t>cV|s-A5173ePcNai0*uvbUt9blb,r7bksozEa8bFa*znBtHXTPa88s1E\\\"\\\",2):f(\\\"\\\"};w7Vtw,Mm*GEEa*FnsizPaVakbb82XwVgbXa6*88O+Aah=VqUaq0N5;2X-fb7lwF?wONx\\\"\\\",2):f(\\\"\\\"}6qQa3J2SBS*X,blw3w2bD>cVIgbFY8g1ubhm4eX,-qG3Wov=UHdbwvKI.b,\\\"\\\",2):f(\\\"\\\"}FaWaET\\\"\\\",2):f(\\\"\\\"}b95Xaf|+yKAtb|7U0A6t>Ra|pEayq8sG:,bxMZa*JL?Rrcb36Qa<aP*+b\\\"\\\",2):f(\\\"\\\"}beQTQAaqXBy=j7cndF<KfdtZ|tbV0y|+b7XnJ|bki><8@UszcCpDPf2P2+b3yFa=rO,2rCpvtGa>H27wuH>HqkiV.0A/ymbe5+bKW?wRzlr>a/u<Rj6-XTtXu9bL6.b,\\\"\\\",2):f(\\\"\\\"}-iWaiss=Zps=9S5b;qNZAq**mbhEYSo\\\"\\\",2):f(\\\"\\\"{9uzpn*l*VxX1:50Rjy,2<t\\\"\\\",2):f(\\\"\\\"{b0v\\\"\\\",2):f(\\\"\\\"}bGYgbqF\\\"\\\",2):f(\\\"\\\"}AqT4DTlrTm"));
$write("%s",("biby7zwc3byrTEaGs971bT2RZtUI26rx:^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3gcaTl^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3c#avydbwFON+beY9b=<Yu-d4<A+RD5b@x?9eY2OXDavzb2Bqx@SIg28\\\"\\\",2):f(\\\"\\\"{z0p;=aeb218VYELx?+;5\\\"\\\",2):f(\\\"\\\"}bxFLDzbbb2bBABf138b7FEaOF.WJ6/5PtQa0q4:/AcxtZVR0tRNzYmQ?v0Vnnfw*1lFPs@wohXarLPN9\\\"\\\",2):f(\\\"\\\"{z@Aaf;\\\"\\\",2):f(\\\"\\\"{pVH?*KY?avb4xO=VHGr@QrghbE+Rm.bTahvdluCvbTaRm*bALvbuBegD"));
$write("%s",("vu/xb3YhYe\\\"\\\",2):f(\\\"\\\"}@,\\\"\\\",2):f(\\\"\\\"{u>\\\"\\\",2):f(\\\"\\\"}=a4b0OEtbbUHBatbVNabx@S4B0O|mLv\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{wgpr.VKwblbCatns=gbWC0bd5Lxlb8b7,dYZas\\\"\\\",2):f(\\\"\\\"}8b9Wm*0rlb-\\\"\\\",2):f(\\\"\\\"}vsp|wAzSU<xUAaw=/sW+3b,zfbvbtHlw=o8C\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{y\\\"\\\",2):f(\\\"\\\"{.P|PHBhxIvuy\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{w15bQuwJabRm6bHz\\\"\\\",2):f(\\\"\\\"{HGsl<O=+wLqpu5\\\"\\\",2):f(\\\"\\\"}kK=\\\"\\\",2):f(\\\"\\\"{g156dsb+p3y|zL|Veb/bVVvtStQ\\\"\\\",2):f(\\\"\\\"{Kp\\\"\\\",2):f(\\\"\\\"}bswL\\\"\\\",2):f(\\\"\\\"}AVzITy*JNCAaCpZo\\\"\\\",2):f(\\\"\\\"}bYE*2>\\\"\\\",2):f(\\\"\\\"}L>KK3bU;DEB.=1KHgbtI9bepnP,Pabyb9r*zNCxhXaVKdr4bms@a,Az|hr5=Cs3sLU+5ub<aGiyjDi>aCp?+GE+deMNrubOVq?UaU>Fa6n3bG:<aVxMO5bCO6bEaq+dLTaTB.bt:;7CE.s.wQycwk?-Qi?P15OBbr0=Sdb9\\\"\\\",2):f(\\\"\\\"}P,Kt-2yb*V|VIGyhb+oMYS7b.s2sSCgbv\\\"\\\",2):f(\\\"\\\"{5byb"));
$write("%s",(",bib4?YEJD|blbdr.bCr?DZamR0b*SCpQ/|+M=-,kb58eq0Fu.GaS/.b:wjb+4y76svIgN;JzbAa\\\"\\\",2):f(\\\"\\\"{bxbDabv>TevUa2b,bQDRaO3PvA16,8j|OkTw-H2eyt,0yTyhVjbZa|9rrZEL-ZaXaAnW|o*2O\\\"\\\",2):f(\\\"\\\"}LP61bvbohj+8wRa96/u=,bqCpOrKx6rL-Qs6-7GJDzbSOt/cQPr71KvOa6-SaOh2Sl>lb\\\"\\\",2):f(\\\"\\\"{wZFYEbuS5+bYB9bKsub*+?aH,\\\"\\\",2):f(\\\"\\\"{kp-vAo4xS.+81P,2b|b:ua;R02>+<\\\"\\\",2):f(\\\"\\\"}bZab*-lGEub?3BA7gC.?ar3R\\\"\\\",2):f(\\\"\\\"}a*8bDaCp>z=wZav7IM5b,PdrW+y,3bfpRa2r8TZ8/zBa5bj1FaTvbvybwb=aQoab95wbcsi+@?\\\"\\\",2):f(\\\"\\\"{b@4VaIq,r?+pCdb+HF-u4dqkbwb1bl\\\"\\\",2):f(\\\"\\\"}x9F4p<Kv2yvzl+0CG,ryepeDCcWa?a3bYqGOJ|Y3gMCQ/4-8@amptbbvK=BvB0bb7q|b8PH|\\\"\\\",2):f(\\\"\\\"}zUa<kAz\\\"\\\",2):f(\\\"\\\"}LNafbBSWq2RWzNa=,\\\"\\\",2):f(\\\"\\\"}PebOa<.o\\\"\\\",2):f(\\\"\\\"{wb.SNCrsRa3b-It*U8WKGaY*Eakb=aUap\\\"\\\",2):f(\\\"\\\"{FkDa-b0\\\"\\\",2):f(\\\"\\\"{*kW<4I/6,Q\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"}skiluORrxSa0\\\"\\\",2):f(\\\"\\\"{6b,C5=X*a7Xa-b=uCs>xcLex2sA06b6bIFe;@RSjTak1OaD2-BKMv\\\"\\\",2):f(\\\"\\\"}j+Z5|mls\\\"\\\",2):f(\\\"\\\"}Lo\\\"\\\",2):f(\\\"\\\"{buPj0bPrfPxbGL-ulbj+0F|+KrAL2O-+O-0RfbSaK?\\\"\\\",2):f(\\\"\\\"{6kb;JUpfby|/trv;t2.g5IG=x-l9yI;:zPa=aWaPaH6ubjRxq5bYAFawbsQ>|xbh;,P4bizVxbbwJtb4=ybkiwI;@|sfbG??2?=ybKvy*Zyq+Ua/uv-s6\\\"\\\",2):f(\\\"\\\"}zbp|/*b3bp\\\"\\\",2):f(\\\"\\\"{zbNaos9x2PCj\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}4w*z\\\"\\\",2):f(\\\"\\\"{K4:Szu<tnQa-i3Fywo4\\\"\\\",2):f(\\\"\\\"}C4M4O,bQjXarx=aosFadb4bMH>3vbk*C.|dC.+cX\\\"\\\",2):f(\\\"\\\"{ubuItbB<MCSrEatsdbRq8blbMOKv:0G>*bNai8PuM4cbVaf*\\\"\\\",2):f(\\\"\\\"{bSag6i+cuHuE++qVvN?9bkb-\\\"\\\",2):f(\\\"\\\"}5F\\\"\\\",2):f(\\\"\\\"}bwbb>>|1lU+wbtx,ufbjbvs*qtb4bbbfuK\\\"\\\",2):f(\\\"\\\"}V:4bS=Za0bQ6PaTagru*KNns,seODa\\\"\\\",2):f(\\\"\\\"{bax?NvbNsZO4b-b>pkpipeDk\\\"\\\",2):f(\\\"\\\"}"));
$write("%s",("bpetV1VoTo96fb<a8bdNH;EIRzBz1bCaz|E+:\\\"\\\",2):f(\\\"\\\"{kp7I5=<0itG+H+\\\"\\\",2):f(\\\"\\\"}bitO+\\\"\\\",2):f(\\\"\\\"}yGs*yEikvLq@4\\\"\\\",2):f(\\\"\\\"{M4>=qL\\\"\\\",2):f(\\\"\\\"{<:VvnqI*j?4KC10bAM7b9tAa\\\"\\\",2):f(\\\"\\\"}b|;4bUiJuFa6x/xBMubJ?H?e+gbUsD2vb-tzp0?t\\\"\\\",2):f(\\\"\\\"}Rabzu4BaFkOaTa9bBvL?h8n9bb/uS5E80bj6xbZalbq1Ca\\\"\\\",2):f(\\\"\\\"{b*bYa<+Aa\\\"\\\",2):f(\\\"\\\"}A2b:zx125d57xvyRaBaR49bmI\\\"\\\",2):f(\\\"\\\"{vv:BqI2<\\\"\\\",2):f(\\\"\\\"}a\\\"\\\",2):f(\\\"\\\"{Ns4>-ze;4b@>6n2bDtXC4<4x1b>FEaXaU6NaIpi6-iF+ubL9G.CwG|yd25nvf.XsWyv<59v<dbv,uuOa3<4:Cw6bxy@aUaWaSaJr0|9bRG4babv4t49wlb\\\"\\\",2):f(\\\"\\\"}K-buuZa7yZ0xFcK\\\"\\\",2):f(\\\"\\\"}bXaUwepdLkbd@H/=q7b\\\"\\\",2):f(\\\"\\\"}GS<5I,6?8*6t6abN?\\\"\\\",2):f(\\\"\\\"{J.b=awFr40bE,Oj2t>alMzbh\\\"\\\",2):f(\\\"\\\"}mb8vu;Sa0bh8BlRapH@aQa+dGgizKxuby;Hp8bTwt5gF0@.bj:hb1bnrtKNaEaP<N<-*GaGx2b<0R5+.hb?aqs0.t"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{Wa\\\"\\\",2):f(\\\"\\\"{DbbWaJv0bjbgKubibK5ib:KD3y7R4c:zbr;:1R>Eav6Mv-+tsCp6b.9\\\"\\\",2):f(\\\"\\\"{bNa=pAxfERa8?85/ber\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"*p=aib3b0bFajbUa0.1zjJdbtb9b;\\\"\\\",2):f(\\\"\\\"{bpUx=1O7wbgbLweJr.F0bkm;Fz>albj>Bagbh<ab3b;595B0590HVx|pMCZaH+4b,\\\"\\\",2):f(\\\"\\\"}4bu\\\"\\\",2):f(\\\"\\\"{Eaxb;9\\\"\\\",2):f(\\\"\\\"}G1IguQaK=I==awbKAo?mbP|abWqk9c+-bC.Tuw95b=5Oa?a9pvb4:h-n+jIOa=aFa/y5\\\"\\\",2):f(\\\"\\\"}i65bcbA1N4S?oJZH@aZ|cbrgxdWaYaH5Zauqy;H?bISa:j1H/Hqi6b7HI>J>\\\"\\\",2):f(\\\"\\\"{9aIRaj=E6/4Ya*bk*@alJV\\\"\\\",2):f(\\\"\\\"{ab=59G,b+cTa1bE69bFaCaUqQaj7SoRaFaoJCqjbhJH@G|7b7HDDVaQa@a\\\"\\\",2):f(\\\"\\\"{bn/wbzbo\\\"\\\",2):f(\\\"\\\"{-bz-3hCpLvMz@>:IVa1xNqe;twRm\\\"\\\",2):f(\\\"\\\"}b/b07bji;4v..IvYaebWalF@a7l.*=aLEzqAxQG<a>ajz?>F8@hgb-2gGKxp|16@8G*\\\"\\\",2):f(\\\"\\\"{C\\\"\\\",2):f(\\\"\\\"}G7bJ76DVaVaM?1@Raxb\\\"\\\",2):f(\\\""));
$write("%s",("\\\"}0cb*bmEGaH36bFa?.5b.q5=x5m3db*qqumbj6db:zF-xb9b8bRayb@a7.<a2Hvb.bAa3q:9Da,bRtzb3udbSa:s0\\\"\\\",2):f(\\\"\\\"{9Gqwwxab\\\"\\\",2):f(\\\"\\\"{2lrE6*swbT/.H\\\"\\\",2):f(\\\"\\\"}HYFtbB2r;Baeb6|v-cbmbhBybNaCpFa<a7bPaDqGoR4mbO-I>6sBaCG<aVa4CJvzb<aOacb1bvBX\\\"\\\",2):f(\\\"\\\"{?>.bzbebybC\\\"\\\",2):f(\\\"\\\"}Aa8bzb-.7CWygb,uz57\\\"\\\",2):f(\\\"\\\"{+bFGwbCBzc6+Ya|,MvkbwyBaOa@ay;ub?@qihb7CT26,xr7zCj7p+c,bX,xbs15b7l.hQqU|wC9\\\"\\\",2):f(\\\"\\\"{hb<.wb7/4a\\\"\\\",2):f(\\\"\\\"{Glq.EOaE6O\\\"\\\",2):f(\\\"\\\"}E\\\"\\\",2):f(\\\"\\\"}??+5So=A56v6?|jb=a;tibCwef,b\\\"\\\",2):f(\\\"\\\"{pcbIghw\\\"\\\",2):f(\\\"\\\"{ba?/z>aDaRa36AuQ\\\"\\\",2):f(\\\"\\\"}dboh5sK/FadsDvtvK=T1,qbp1bz9Afdc/p@DogZyebHC\\\"\\\",2):f(\\\"\\\"}uzbW;yjPamb|/q:TaiDDa*\\\"\\\",2):f(\\\"\\\"{cbm*k*\\\"\\\",2):f(\\\"\\\"}bRaM4W:y9w9Cau9J4qud?Is0btb?xmb2ymbcjhblbz3\\\"\\\",2):f(\\\"\\\"}b.bXaR1<3=,I/mb8ba*\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"{yWaCpCqeb0b9f@uG:+88gOxhv-t4>:|OAd|Fa5bo759O,Cpz;Ba-b\\\"\\\",2):f(\\\"\\\"}b?0X*tEL\\\"\\\",2):f(\\\"\\\"{9sHv,xyD07W3?|/+VwN5VaG,R*ns4vvk,ED*yCBa19guX*TA\\\"\\\",2):f(\\\"\\\"}b1>m*@a4>Op0bwbWyu;Oy+:E.5sXo3b9fd?fkBaAa*bS=r/lwki8tG:ubF+hr9>7bM8ub0b5@07.dU5fbMzZaXua?4wzb2*Da=pNa-tcbybA+9w7>gbffwDKAQuNaSvfbdb:6qsFx:5G:7|Sa1bVayb1bUaDaAa9bZambxbkbDpT\\\"\\\",2):f(\\\"\\\"{g-z5+zebd:b:;1Y9,x-\\\"\\\",2):f(\\\"\\\"}ib/tUa28*,=af.ib17Sa|b<a/xzd>azpX@7b*/TaZad\\\"\\\",2):f(\\\"\\\"{Uz8bFBl\\\"\\\",2):f(\\\"\\\"};w+qA=-ro7j72**b.bGa9B312*H?g9+bhbnw;1-b3yDahy>4bbo\\\"\\\",2):f(\\\"\\\"{,b92cpp|h?BytA*krARa-bGa;<\\\"\\\",2):f(\\\"\\\"{u1yDao\\\"\\\",2):f(\\\"\\\"{9b,u|2Va|+2b*b7\\\"\\\",2):f(\\\"\\\"{g+ZpFx/4xbAzxbB\\\"\\\",2):f(\\\"\\\"}Sl2bJ2-=BzNa.bTlSxAr?-Bw7bcsBa/bLyI8Say|Ya3\\\"\\\",2):f(\\\"\\\"{|+cbO>Oag+n,B\\\"\\\",2):f(\\\"\\\"};+ixjpcmV8wbBqabEr2bPaDlA5c*ubFs"));
$write("%s",("/bubFa\\\"\\\",2):f(\\\"\\\"{b<aV:CqY0w11bKq<ak9cshu5b>.a94b,bfBfsMwR1/:zbb+Os++\\\"\\\",2):f(\\\"\\\"{2e+Uwg2Y7kbD9Wreb?\\\"\\\",2):f(\\\"\\\"{d*,>9ukwGr8b5b1bAzZaBazbbkO-1\\\"\\\",2):f(\\\"\\\"}bz=9+p@aTasuW2t>\\\"\\\",2):f(\\\"\\\"{bJ|?-8gSx5bb/=acbCps=53RmEavbnwbclY2bmb6xtbypvb?nHzcwm-V<*kT<\\\"\\\",2):f(\\\"\\\"{kR<zb+b5z,po9Za|pbcWaAaU?;qjbebJt=o+z\\\"\\\",2):f(\\\"\\\"{j/bFa\\\"\\\",2):f(\\\"\\\"}bu4GqC\\\"\\\",2):f(\\\"\\\"}ns|8Xa8xCqk@8/jv>@tbhbjb0b8bwb*\\\"\\\",2):f(\\\"\\\"{fbu,h/Pa@ayb@4kiGtUanvSaebe@8bm@ArBaEayb81=5Rar<mzSzY.5<?+UaubebE+Arg6T6*b3qo7@a9sEa/bc|4bk0=aSzRaU?b+zbF;PaxbdbF>81yxeb2bFvQa1b*1A5J7<kgb9b-bkvfb8b-b8bazB?zj>i?-BaubTqdz3b7buxOyQxLt7qB\\\"\\\",2):f(\\\"\\\"}7bQacbSaXa<a>|+5|b90Xa9zr99sTatbaizpCjVi2uLrU0Yavb.9QxZanqZvg?N:lt+6j4<t12?\\\"\\\",2):f(\\\"\\\"{CadbxrxbS+Qa\\\"\\\",2):f(\\\"\\\"{d|b5:?|Xay;u4Wa2s8bdbubSaJv:w|;1b<s*|5"));
$write("%s",("bb;j>Xa>a72I4ybjb-q5b3b\\\"\\\",2):f(\\\"\\\"}bslR5eb5b6bXa.xS1\\\"\\\",2):f(\\\"\\\"{b|bRalv7gEaz0;.9bpsp\\\"\\\",2):f(\\\"\\\"{abhpabib*bXakiw5,xnn?qWaF+8b2\\\"\\\",2):f(\\\"\\\"{kze/xb8bdyJdCpsuquOahb|sabU\\\"\\\",2):f(\\\"\\\"}Ux6bUz|bEtNaybX+=7wb\\\"\\\",2):f(\\\"\\\"}bdbTv2r/sLqBzLqlw6x?w1bhpm,s+f+H2\\\"\\\",2):f(\\\"\\\"{3Dar.ub>a\\\"\\\",2):f(\\\"\\\"{bhbFa9\\\"\\\",2):f(\\\"\\\"{xb7bkb.br=0b>||/B\\\"\\\",2):f(\\\"\\\"}<.xyI8A,F-|b+sMrxb\\\"\\\",2):f(\\\"\\\"{bgbefQpB0jb?vxpFaCqFq=a\\\"\\\",2):f(\\\"\\\"{27/\\\"\\\",2):f(\\\"\\\"}<Sa@<ki?17b\\\"\\\",2):f(\\\"\\\"{kB*06\\\"\\\",2):f(\\\"\\\"{kE*o4O:VaG|mb/*t<O+Gog.h..b2\\\"\\\",2):f(\\\"\\\"}Ean/AaSjub>|vbCp;uubkiw/mbVaCpguu-Ca7blb+.,rkb81JrSnf.XambY-48Jrt<WaRa<.lbIqSambUa\\\"\\\",2):f(\\\"\\\"{.zjUiRaHp/b,q4b+bNa0\\\"\\\",2):f(\\\"\\\"{g1=wyqe/TaLq4wA,kbSzg4jb|\\\"\\\",2):f(\\\"\\\"{ab1\\\"\\\",2):f(\\\"\\\"{6b=q*.t,fgg;e;1w3bkb=kYa+pLxk;O-w|0byyx|j3eqC\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"}Pa9b-.9ft*G,QaP|frNhK\\\"\\\",2):f(\\\"\\\"{?fx9Nav:***zS+Bawm3bXaTarj\\\"\\\",2):f(\\\"\\\"}smb90dyOaO+3bKzIz3bKxC9YaVa>aQalb\\\"\\\",2):f(\\\"\\\"}b5bibsv4bS*F2\\\"\\\",2):f(\\\"\\\"}9\\\"\\\",2):f(\\\"\\\"{9Ya8uy75uHnqsp|M:?y=8FxN|Pa+ynjbbib04SokvI8\\\"\\\",2):f(\\\"\\\"}/?ah:z9Dr\\\"\\\",2):f(\\\"\\\"}bD24vx3ak=p6bVaBah:+bI8-h,bypvtPadb6z1x,b3q/bRa?aex\\\"\\\",2):f(\\\"\\\"}bjbcrRaJ/ybHpT6lb?a4\\\"\\\",2):f(\\\"\\\"{=27bm\\\"\\\",2):f(\\\"\\\"{/bbbc:pr3bTatxPadzUaEajuA\\\"\\\",2):f(\\\"\\\"{I49z95ib\\\"\\\",2):f(\\\"\\\"}.*bbbbxUaMvU-l/Twx-OoNpWribVadbxbv0lp*bOxt\\\"\\\",2):f(\\\"\\\"{FaV\\\"\\\",2):f(\\\"\\\"}L6N4jzgbQag-TiXj.bVaxr@\\\"\\\",2):f(\\\"\\\"}4bN*R*nvUa8b|bub6bDaQa2xkbAa4bv-;*PrWa9bC+Ta\\\"\\\",2):f(\\\"\\\"}bPaScTaOa@0p1R8YaYg6b|bZaC\\\"\\\",2):f(\\\"\\\"}W+lbBakbJyvbtwUtfbZafbCpBak+Za|+?+jbfb18W+nq-6O1m4M1k4-b7/58X5Fa?,.+8b3b\\\"\\\",2):f(\\\"\\\"{bfbCa3bzjTaSa8/c"));
$write("%s",("bz5Dzps\\\"\\\",2):f(\\\"\\\"}6Xa\\\"\\\",2):f(\\\"\\\"{6UqVaDa|7v6M6jy>a.+V1PaW7U7@5MttbwbwxQ\\\"\\\",2):f(\\\"\\\"{Y3Rm25tuz2y7NaQ7cb>a|bgb1b1l<a46dp176pE7Ralbvbu4+zCpvb:whbN*=,=afbFa3blbjbQxabp1xba7Fahb-iu,5bCaQahbtpHjibv.x6tbN6L60bolm7>an+VwT2wb:wvbVags46dr*b@a.,fbTakbu,ysjyhb,bL\\\"\\\",2):f(\\\"\\\"}6b@aDacbFaxbQxG-vbDaw6fgabgbgb4bXzhbybJyhb:p\\\"\\\",2):f(\\\"\\\"{v-2Huq\\\"\\\",2):f(\\\"\\\"}3p.b364bLqQaibkpGqGrcbtbjbcws|n4p|l4o4CyN1J1O-Nx>a+|xx5bb4.bv|/*wb*bwswvLy.btwSsWa|b@aBaabTvD+B+Sjwx\\\"\\\",2):f(\\\"\\\"{bdb+b3bF-:zGskb7btb@-zscbEa20PaRawvM|5z\\\"\\\",2):f(\\\"\\\"{yXaecAaxbL\\\"\\\",2):f(\\\"\\\"{gbRaYqE+Sa\\\"\\\",2):f(\\\"\\\"{bZaQa9bQa|x=,HrfbfgYab,zbCaTa=,rp*bZ2fbz|/tAaPwCpDaJ4dqabAaH,xbYm-bxut4Ra.-sl\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}JxzbXaYwQaeb\\\"\\\",2):f(\\\"\\\"{bQaDaEz43tbrvHzI4\\\"\\\",2):f(\\\"\\\"{pzbR\\\"\\\",2):f(\\\"\\\"{dbhb4b"));
$write("%s",("CaAa82bbmb0zh.=aR+6+E.>|@a3bCp2bQa/t/z93>\\\"\\\",2):f(\\\"\\\"}Fa1x-dybr4i4njg.,bkbQadb8bTalb.bp3@i\\\"\\\",2):f(\\\"\\\"}b*.f/cj*b/b4b8u*bcwL1q-D/cwB/K10b*3+bkb\\\"\\\",2):f(\\\"\\\"},Y0ai>i8bVa7b>aUaUaibFq3s9\\\"\\\",2):f(\\\"\\\"}+bAxabRtdpdcTq1bebHx4svb+v.bSaVobcqugk3\\\"\\\",2):f(\\\"\\\"{|bHscb2bLxgbLrTaX2xb?aFgibCa>|6bUalbScqu2bbq6b2bcbBaxbvbGoFg@2GaC,ibubybw\\\"\\\",2):f(\\\"\\\"}Baiuky7bohCqMqbb82cbfb/bfbbbTaWa0b>acb\\\"\\\",2):f(\\\"\\\"{b@2|-bcQai|X/|bTl8b,bfb|b.s3b2uQa9scb5w1bQa1sjuWajb0w-bAa@aGagyVwnwolZahbtb@aFaYa3bybPa+b@akb0r=aXqU+J|wbo\\\"\\\",2):f(\\\"\\\"{ace\\\"\\\",2):f(\\\"\\\"}<aJsPaQ/Lqo\\\"\\\",2):f(\\\"\\\"{yxMstbPa>|fxXuCaabV1kbwzAsyy=aB1+bab?asqE/qtC/n-dw@/2bLsz,juAujrt-Ua|f/bG,PaF0Na7zYa?a|b2bdb8zvbjsBaYa:uj1bbW|Ssz*e|vbY\\\"\\\",2):f(\\\"\\\"{G0fbEv1b5b/b7b+q?aNa@pkbgbM|Ip-xM04blbYakwWappwb\\\"\\\",2):f(\\\"\\\"{0B\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{,qab0bXa=avblb,bubWxXaJhwy0ptsFaG0zsVa8wVsUaeb-\\\"\\\",2):f(\\\"\\\"}7\\\"\\\",2):f(\\\"\\\"{0pNa0b@atb,xCaDaD-abtbL\\\"\\\",2):f(\\\"\\\"{CaKzI-G-E-a.B-0b@-VzFg<-:-ubPa7gfx\\\"\\\",2):f(\\\"\\\"{bmbLqHs1b>a5w7vm0hbG,hcwv|bS|gbg0Pa>a3-WqX.QaU/OaU/SaU/NaU/w.R-kiNt\\\"\\\",2):f(\\\"\\\"{tRas-LtEa1bHjbyOaWaXab*9mp|H*nqawyio-Xa0b..z/c.7b/bVaUa+bcbp/u/s/Ra+.=uJr?a1bBr4bvb0b4.EaO+;*@aL.=aSadbNa@a+eAaVarv7bc.r.gbdbYmlbeb?aaibbYmc.jvdbCp>anvb.1h1bM|L-dbDadl0-ib4.=aVaw./bOaSa8b*bSafv+b?aX-mbXaUaAqu-.b@ac.=a\\\"\\\",2):f(\\\"\\\"{bOaa*BalbRa8b1hRa>aEaAaSa6b+bY->aSaub+bakAampFaY-3bmb|wgz?q@aWaWaTa<af-RaAaeb@aSa?aSaVaSaAaOaNaDt|,abM|kbmbKzYaFsabCaxbLtAaYuibqu*bAauxirFiibebCaPa3bParz0u6bxb>a+b9|?a\\\"\\\",2):f(\\\"\\\"{bFaau+bSo6b*bkbSaybXalbVa?af-yiF*Eyl-mtqoA**b*uquibEa.bGpvbybgbkbBaXaSa4xS+Di1b7bqw>aPa/b@ax+"));
$write("%s",("*wCaq+1bhbCpk+hbx+:rNa?ak+Dae+7b3h,dgu4umb>aFahc9uS+lb@aXa\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{Fa/pfbybQaSatb+blb3bq\\\"\\\",2):f(\\\"\\\"}.bOamb/bLtmubb>a-bXa?aWabu.bkxbbjbXs4uW*gb\\\"\\\",2):f(\\\"\\\"{bfwSa@hBaCpkbLxzpSa.bSjKsgbyh-d:+8+\\\"\\\",2):f(\\\"\\\"{u+|>aK\\\"\\\",2):f(\\\"\\\"}4bYaDaubWatbyy\\\"\\\",2):f(\\\"\\\"{bnj:t,ber:uzb9yRacb+|vuzb@a++ZqkbNazbAzPa1bYqNar+?hTlki|r*bjbOazbbyCprzO\\\"\\\",2):f(\\\"\\\"}0b1lGa>*lb-b/u@a-bfbi\\\"\\\",2):f(\\\"\\\"}1bPa*qkimmibzbax4btbdq0b/bCatb0bC|Jwbb9mcwiovkC*@y\\\"\\\",2):f(\\\"\\\"{in|o|r|Caki:*<a+bCp0b\\\"\\\",2):f(\\\"\\\"{b5bkjPa7qWq:x|bMhYrWacbz*nv?a0b+bPaFakbtbSawbjbPa0bhmTub\\\"\\\",2):f(\\\"\\\"}wbcbbb\\\"\\\",2):f(\\\"\\\"}babYai\\\"\\\",2):f(\\\"\\\"}kb+jsu2b9rVa0bOaXa4b\\\"\\\",2):f(\\\"\\\"{bPaibAawbIoVo0bUa-bOa?sF\\\"\\\",2):f(\\\"\\\"{vbWa:s\\\"\\\",2):f(\\\"\\\"{zkb|\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{j4bfbQaBaTa+bQa4bT"));
$write("%s",("i/b|bns,bQuHpfwcb\\\"\\\",2):f(\\\"\\\"{xyxQaTa;vnxdqibbbLj?a6bubkb\\\"\\\",2):f(\\\"\\\"}v?v2bYaNa\\\"\\\",2):f(\\\"\\\"{b6bvbXaZaPatb|bab|bdpvb<aF\\\"\\\",2):f(\\\"\\\"{8bipZaYwLq*bc|Cp1|Vz*b+b,bAujb:pVrubZaibSa5s-dBaUaTaUaMuC|A|Ea\\\"\\\",2):f(\\\"\\\"{b?v,xQa8bYay|kw?aub.b,bbbabEiQuFaOa/bjp-tXuibjbXa,rQuPofbebtbAaPz*bnq|km|IbFy>yyi<yNy?w7bSaYwq\\\"\\\",2):f(\\\"\\\"{o\\\"\\\",2):f(\\\"\\\"{m\\\"\\\",2):f(\\\"\\\"{WazbUa3v6bwbNa4b@afs4pNa3b8bgbBar\\\"\\\",2):f(\\\"\\\"{OsUahvWyebr2=lCaFa;\\\"\\\",2):f(\\\"\\\"{=\\\"\\\",2):f(\\\"\\\"{PahbBaJtDatbNa9bUaLq.babNa<tPa-bdbVaFa-b3z.dxyQoZxybervbUa5bVaPwef=abbQa-bFaQxkbOaibab*bQa5vrxYatzrz=kAa*z.x|b|bVzhsAatbbbTvubdbsxXaGu?z3b+bdbabTa/b=a/bmbab7bZaUaOatcmbQybj/bSabbwbPaXaRakbhbhbcbAa5b6y+b>aababbbrzDampsuYxzbhbIp9v.bDaldwbYa|bVaXaDa/bAaAa<a\\\"\\\",2):f(\\\"\\\"}bLxfbVrtbVa8bMqhjOa5v/yTaetAaTaQxEaYaYumb"));
$write("%s",("VxybmbevyiDystAypqpt=yntcwrqvkbwUa/b\\\"\\\",2):f(\\\"\\\"{bIhLxyy7bdp\\\"\\\",2):f(\\\"\\\"}bNa1bWx7brrOpljjbibdbyyibTi8bWa1bcb3bPrGa6vExgrCpmbivduVx\\\"\\\",2):f(\\\"\\\"}b?nkiOvzsab\\\"\\\",2):f(\\\"\\\"}b<a?aabuqQuouubgbib=a*bcb8b/bXaeb4rYaabEa@ukiBp6b@xAxCp-u,b<tRaXaNaWqxbXaibtbOa1b8bmbCa-b*bVvbblbibTaqpXa4e*b=aYaRaDaUatbcb|b4bhbVtHg:vEa0b\\\"\\\",2):f(\\\"\\\"{w\\\"\\\",2):f(\\\"\\\"}bcbgb5bEadb1bbb\\\"\\\",2):f(\\\"\\\"{bub9bmbcbXavb5bvbwbebhmYaFa,b\\\"\\\",2):f(\\\"\\\"}rwbZaAnVaxbLqzbmp,bpskbeb@iyw0b@gFamnkbcb5bNaXaLrib>aubSj,bZa6b.bfr\\\"\\\",2):f(\\\"\\\"{bCphbabcb7bXaQakbEaLvYa.bWars*bTamjOaDvtb\\\"\\\",2):f(\\\"\\\"{b/bcb6bmbBa9m4attYvlonqktgbOrYa=a3b5bStQtOt-bEaebQa|b/bUacbCa\\\"\\\",2):f(\\\"\\\"}bYaQa\\\"\\\",2):f(\\\"\\\"}b+bKugb*bCssv1b9bxbAajbkiar\\\"\\\",2):f(\\\"\\\"{bAazbKu1bfb,b6tLrksdb4uybUkEalb9pvuCphp4bWaUa>a5bZa3bCaXa\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{b8bOa=pzbSa=adb:jIu*bPqeb\\\"\\\",2):f(\\\"\\\"}bEatbLuAa>a@p-dgbmbmbhbgbubbb.blbSacbdqvpybybOa2b1b:tOaEaep5bYacb4bgbdq,b=a1bwb@aOa3bvq6bkbmh/b-bRaUajbwbyb8pmbgb+b8b0bdb,bPalbCp\\\"\\\",2):f(\\\"\\\"{bEidb3bOaAaFa1bSaabQa?axt4bAais,b6bTaab4beb|bCp?a*b7bFaibHqCpyblbTagbZbBrWaKoFa3s1s5bwbCaCpib7bibQaKrkbWa*bFaeb3b,bWaCaebvb\\\"\\\",2):f(\\\"\\\"{lwbTa\\\"\\\",2):f(\\\"\\\"{bys?azbyirtjqotoo,mqqmqnq<mgqBrjbssqsoslb9bksisgsGaes@a/bPaWaQc<avbQawbwb7bNa/blblb+bXaabwbmbubvb\\\"\\\",2):f(\\\"\\\"{b7b,byb/b<aib-pWaEaCpfhubCp\\\"\\\",2):f(\\\"\\\"}blb6bdbwb2b0bCahb>aRaablb\\\"\\\",2):f(\\\"\\\"{b-bybfg>aebjbTaYa,b-b\\\"\\\",2):f(\\\"\\\"{b1bkb9b.b?aebgb2bUaki1rRa0bJqTacblb>aNaYa0b=aDadblb5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaSaCaub\\\"\\\",2):f(\\\"\\\"{p9bzbjbRazb2bVaTq,rNoCp.bCaXq7bfb-b3bUaCp7bVatb.b7b2bfrdrbr*b3gUavb@a0q/p\\\"\\\",2):f(\\\"\\\"{bCq"));
$write("%s",("Uqdbyb\\\"\\\",2):f(\\\"\\\"}bkbdbkb4bjb-b7bdb0bPa,bOaxbCp,blbUaQa>aib,bebVajb,b0b0bWaBaFa+bSaEa4bUa|b\\\"\\\",2):f(\\\"\\\"{bebmb3bDa-pmbTpzb=aTaNp*bBambPaKojbFaPaCambFa>aTafbibOaCajbhb6bBa9bPa|bAa-pnqko\\\"\\\",2):f(\\\"\\\"{ihq:mkqmoyiiq/mpozknomb0bcbOhjbkbPa4b=phbNaBaDamb4bBaibwbhbvbkbvb3hZakbibnhlbGa5p+bfbwb5bXabbCa|pyb0bfbYakiqb4bDaYadbvbzbnh|bbb5beb|pjbcbwbWaNaDa9btbtbDavbhbPaEa+dXazbcb.b-beblbzb,bNa7bvbCaEahb<aCabb*b8hQaub*bWaQagbSa,bEa7b6bAaEaUm>ofn*owouoXf*o*n?aSg4o;a2n\\\"\\\",2):f(\\\"\\\"}nuo\\\"\\\",2):f(\\\"\\\"}oQm.o-b*o1nCa/nWnwbic8aZnEnFmxoEaQmFntn-a8npnnn9m\\\"\\\",2):f(\\\"\\\"{ijo;mho9a9m*k*k-m9m/b\\\"\\\",2):f(\\\"\\\"{f-a;hub@h|eQnIn<nMnDm9aEaOa>mvnGm/nVmzn2i:a>n=aAa/n;nCafnwn-n@a<a-b2n6nWm2nYmEm.n1nAa:aCa8a+n>aXmPmenZmKmhnAa0lWm|eqnzbHmbnImSmBaEmOmMm*bvbtb/b-aJdHd>manRmWmUmSe|eNmTm?aAa-"));
$write("%s",("aDm8aJmHmFa@aEm\\\"\\\",2):f(\\\"\\\"{bCmHaAm9a|eBmxb8a+e-a1beg>mum8arb8aXf9m9mMi+k0m6l@l,k7e,j*jokyi.mvk+myk\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}knm*j6b-a+czbxbubHaqb6aqbEiFiDi5aqbebYi,bAfzb.bKfnbxb\\\"\\\",2):f(\\\"\\\"}ikiZgXgagIkAl2j.kel?a=aLi;dLf7lRi5luh3ltcBa3aPhIgDiwbPf?aRkYkNkBa?aKi6e;hrbTk?a7iQkvhOkDa?a>aKi2b3bGiUfTj8f2i-b:kCa3aKa\\\"\\\",2):f(\\\"\\\"{b;a3gwbccIa3b1bbk,b|b0auh\\\"\\\",2):f(\\\"\\\"}h6hlk1jjkCaKi.bti0kkkMi.jyb3bKk7hDh/k*h-kBaLiMf1i\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{gsbubwbki-a;k9k:a;b6k1b0b-b3aAa3a7b-aki.a:b:b,b?a3j5i5h0jik4axi\\\"\\\",2):f(\\\"\\\"{k\\\"\\\",2):f(\\\"\\\"{kwk3aLiyiuk-fzi-j5e+jmdrjRf7hvhQiOi/j3a;hwb+b-aPcPj/b8b1bPcxb;aUf-b:fZapg|b.b5b-aHj>i3bWfvb|bIgGipgfg3bgf;a<b:b3b-a8bIg,bxb2b2btb;a7hWhPimiNi@aKiIhujxbsjqjabVaTaRaOaHa6eEfOhFfjb-agbebbbcbZaVa-abbVaEf-aZabbebSaHa@g-a3h"));
$write("%s",("hbQabbZa7h*h6iPa4i3a>a3a5anb-aEi/b3b4b.bHa8byb2b2gtbWfxb5b+bYg7h5hliYhWh;d+cKfHa-i-iFaGaji|fld4a.gwi/auh4a-afgdgMaFa=aWh-bYhDhChGa+bJdRh9a/b5a|fCc8g-bPaBaobDhHfMa9aMaIa5axb3b.b4b0bxbzb-btbeg7hkg5hGaMbHg2bzb;azbLfccJa7b?a?auh*hCdYaOaVafbVaibNa=avhvh?a;aSg\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"VaNaUa.guhkgvbpbEa*c7bDaFa?aDa>anbJdubSczbPfIcQgyfwfuf2bsfNd3bHa?e-a-fZf:aIa+c9f:avbldub4bcb-b3ggc0gHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bdgfb/akgzgtbxcRf?a1akg-a6a5bhg>azd:a,cNahgwb.b;b>aagob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a,fPcFf/b:b6aKa6e1b4eIa8btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8"));
$write("%s",("aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,13&X3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)"));
$write("%s",("v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalcz4rfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajm4bdateg@3doa2 kcats timil.v3dga]; V);Q4aC3ecaL[b5aX4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.<5joa(=:s;0=:c=:i;)|4ajaerudecorp/3fqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{.3bianoitcnufR6\\\"\\\",2):f(\\\"\\\"{sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3mja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(ga36(f\\\"\\\",2):f(\\\"\\\"{#j4[j4boa(etirw.z;)tuo.N8aba(67b~auptuOP"));
$write("%s",("IZG.piz.litu.avaj wen=zG4Zka91361(f\\\"\\\",2):f(\\\"\\\"{#tm4[m4c5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/@4[@4cda*6 Q5[p4dea1312^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[w8[$5ofa41310r4[r4c7=[B>[j4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6pma(amirpmi oicy4[(5[j4hma++]371[]591[?6[?6cpani;RQ omtirogla\\\"\\\",2):f(\\\"\\\"{4[\\\"\\\",2):f(\\\"\\\"{4cua;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"})48z3b(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632N4Zsa7218(f\\\"\\\",2):f(\\\"\\\"{#(tnirP.tmfIIcfacnuf;&4[&4bdatmfn4[n4cgaropmi;ILagagakcap~4Zea1304T6dbapD6[r4cba-l4[l4bjatnirp tesY>[ca89&AafantnirK7[ia959(f\\\"\\\",2):f(\\\"\\\"{#fp4[ga^64^\\\"\\\",2):f(\\\"\\\"})74[8awa,s(llAetirW;)(resUtxeT:Paca=:R6[ba1Q6ak8ap4[p4adaS Cn4[vEaca&(z5[z5aba 06[06[06piaRQ margo^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[t4cjaS D : ; R-5[%L[j4[j4o%6[k4aqa. EPYT B C : ; Az4[56[j4[j4nka)*,*(ETIRW/6[J7chaA B : ;s4[s4aba [2cr4[*5dia: ^1^\\\"\\\",4)"));
$write("%s",(":f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohce4B[ka3(f\\\"\\\",2):f(\\\"\\\"{#(stup;Rcdatniy4/ca0153.ea%%%%m4[m4[53ipaparwyyon noitpoz4023[230ca(nVO.ba5FQa\\\"\\\",2):f(\\\"\\\"{aetirwf:oin\\\"\\\",2):f(\\\"\\\"})8(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3c\\\"\\\",2):f(\\\"\\\"{P)ka(f\\\"\\\",2):f(\\\"\\\"{# cnirp/L)l;eja.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[(3rba@~Wa7;alaM dohtem06x*3c|5aV;cpadiov;oidts.dts &Ya;6n+4d\\\"\\\",2):f(\\\"\\\"{3kkaenil-etirw~5dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea"));
$write("%s",("^128^+Ac/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing b"));
$write("%s",("owl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\","));
$write("%s",("9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:Ou"));
$write("%s",("tputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule